`timescale 1ns/1ns
module Q1(input[15:0]inN,inM, input inC, input[2:0]opc, output logic [15:0]outF, output logic zer,neg);
	always @ (inN,inM,inC,opc) begin
		neg = 1'b0;
		zer = 1'b0;
		outF = 16'b0;
		case(opc)
			3'b000: outF = inM + inN + inC;
			3'b001: outF = inM + (inN >>> 1);
			3'b010: outF = inM + 1;
			3'b011: outF = inM + (inM >>> 1);
			3'b100: outF = inM & inN;
			3'b101: outF = inM | inN;
			3'b110: outF = ~inM;
			default: outF = 16'b0;
		endcase
		if(outF[15] == 1)
			neg = 1'b1 ;
		else
			neg = 1'b0;
		if(outF == 16'b0)
			zer = 1'b1 ;
		else
			zer = 1'b0;
	end  
endmodule

module NOT(A, Y);
	input A;
	output Y;
	assign Y = ~A;
endmodule

module NAND(A, B, Y);
	input A, B;
	output Y;
	assign Y = ~(A & B);
endmodule

module NOR(A, B, Y);
	input A, B;
	output Y;
	assign Y = ~(A | B);
endmodule

module DFF(C, D, Q);
	input C, D;
	output reg Q;
	always @(posedge C)
		Q <= D;
endmodule

module Q1_yosys(inN, inM, inC, opc, outF, zer, neg);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  input inC;
  input [15:0] inM;
  input [15:0] inN;
  output neg;
  input [2:0] opc;
  output [15:0] outF;
  output zer;
  NOT _1212_ (
    .A(_1193_),
    .Y(_0928_)
  );
  NOT _1213_ (
    .A(_1194_),
    .Y(_0939_)
  );
  NOT _1214_ (
    .A(_1195_),
    .Y(_0950_)
  );
  NOT _1215_ (
    .A(_0456_),
    .Y(_0961_)
  );
  NOT _1216_ (
    .A(_0463_),
    .Y(_0971_)
  );
  NOT _1217_ (
    .A(_0479_),
    .Y(_0982_)
  );
  NOT _1218_ (
    .A(_0464_),
    .Y(_0993_)
  );
  NOT _1219_ (
    .A(_0480_),
    .Y(_1004_)
  );
  NOT _1220_ (
    .A(_0465_),
    .Y(_1015_)
  );
  NOT _1221_ (
    .A(_0481_),
    .Y(_1025_)
  );
  NOT _1222_ (
    .A(_0482_),
    .Y(_1036_)
  );
  NOT _1223_ (
    .A(_0468_),
    .Y(_1047_)
  );
  NOT _1224_ (
    .A(_0469_),
    .Y(_1058_)
  );
  NOT _1225_ (
    .A(_0470_),
    .Y(_1069_)
  );
  NOT _1226_ (
    .A(_0486_),
    .Y(_1079_)
  );
  NOT _1227_ (
    .A(_0471_),
    .Y(_1090_)
  );
  NOT _1228_ (
    .A(_0457_),
    .Y(_1101_)
  );
  NOT _1229_ (
    .A(_0473_),
    .Y(_1112_)
  );
  NOT _1230_ (
    .A(_0458_),
    .Y(_1122_)
  );
  NOT _1231_ (
    .A(_0460_),
    .Y(_1133_)
  );
  NOT _1232_ (
    .A(_0476_),
    .Y(_1144_)
  );
  NOT _1233_ (
    .A(_0461_),
    .Y(_1154_)
  );
  NOT _1234_ (
    .A(_0462_),
    .Y(_1165_)
  );
  NAND _1235_ (
    .A(_0472_),
    .B(_0456_),
    .Y(_1170_)
  );
  NOT _1236_ (
    .A(_1170_),
    .Y(_1171_)
  );
  NOR _1237_ (
    .A(_0472_),
    .B(_0456_),
    .Y(_1172_)
  );
  NOR _1238_ (
    .A(_1171_),
    .B(_1172_),
    .Y(_1173_)
  );
  NOR _1239_ (
    .A(_0455_),
    .B(_1173_),
    .Y(_1174_)
  );
  NAND _1240_ (
    .A(_0455_),
    .B(_1173_),
    .Y(_1175_)
  );
  NOR _1241_ (
    .A(_1193_),
    .B(_1194_),
    .Y(_1176_)
  );
  NAND _1242_ (
    .A(_0928_),
    .B(_0939_),
    .Y(_1177_)
  );
  NOR _1243_ (
    .A(_1195_),
    .B(_1177_),
    .Y(_1178_)
  );
  NAND _1244_ (
    .A(_0950_),
    .B(_1176_),
    .Y(_1179_)
  );
  NAND _1245_ (
    .A(_1175_),
    .B(_1178_),
    .Y(_1180_)
  );
  NOR _1246_ (
    .A(_1174_),
    .B(_1180_),
    .Y(_1181_)
  );
  NOR _1247_ (
    .A(_0950_),
    .B(_1177_),
    .Y(_1182_)
  );
  NAND _1248_ (
    .A(_1195_),
    .B(_1176_),
    .Y(_1183_)
  );
  NOR _1249_ (
    .A(_1170_),
    .B(_1183_),
    .Y(_1184_)
  );
  NOR _1250_ (
    .A(_1193_),
    .B(_0939_),
    .Y(_1185_)
  );
  NAND _1251_ (
    .A(_0928_),
    .B(_1194_),
    .Y(_1186_)
  );
  NOR _1252_ (
    .A(_0456_),
    .B(_1186_),
    .Y(_1187_)
  );
  NOR _1253_ (
    .A(_1184_),
    .B(_1187_),
    .Y(_1188_)
  );
  NOR _1254_ (
    .A(_0928_),
    .B(_1194_),
    .Y(_1189_)
  );
  NOT _1255_ (
    .A(_1189_),
    .Y(_1190_)
  );
  NAND _1256_ (
    .A(_1195_),
    .B(_1189_),
    .Y(_1191_)
  );
  NOR _1257_ (
    .A(_1172_),
    .B(_1191_),
    .Y(_1192_)
  );
  NAND _1258_ (
    .A(_1193_),
    .B(_1194_),
    .Y(_0489_)
  );
  NOR _1259_ (
    .A(_0928_),
    .B(_1195_),
    .Y(_0490_)
  );
  NOR _1260_ (
    .A(_1195_),
    .B(_0489_),
    .Y(_0491_)
  );
  NAND _1261_ (
    .A(_1194_),
    .B(_0490_),
    .Y(_0492_)
  );
  NOR _1262_ (
    .A(_0456_),
    .B(_0463_),
    .Y(_0493_)
  );
  NAND _1263_ (
    .A(_0456_),
    .B(_0463_),
    .Y(_0494_)
  );
  NOT _1264_ (
    .A(_0494_),
    .Y(_0495_)
  );
  NOR _1265_ (
    .A(_0493_),
    .B(_0495_),
    .Y(_0496_)
  );
  NAND _1266_ (
    .A(_0491_),
    .B(_0496_),
    .Y(_0497_)
  );
  NOR _1267_ (
    .A(_1195_),
    .B(_1190_),
    .Y(_0498_)
  );
  NAND _1268_ (
    .A(_0950_),
    .B(_1189_),
    .Y(_0499_)
  );
  NOR _1269_ (
    .A(_0961_),
    .B(_0982_),
    .Y(_0500_)
  );
  NOR _1270_ (
    .A(_0456_),
    .B(_0479_),
    .Y(_0501_)
  );
  NOR _1271_ (
    .A(_0500_),
    .B(_0501_),
    .Y(_0502_)
  );
  NAND _1272_ (
    .A(_0498_),
    .B(_0502_),
    .Y(_0503_)
  );
  NAND _1273_ (
    .A(_0497_),
    .B(_0503_),
    .Y(_0504_)
  );
  NOR _1274_ (
    .A(_1192_),
    .B(_0504_),
    .Y(_0505_)
  );
  NAND _1275_ (
    .A(_1188_),
    .B(_0505_),
    .Y(_0506_)
  );
  NOR _1276_ (
    .A(_1181_),
    .B(_0506_),
    .Y(_0507_)
  );
  NOT _1277_ (
    .A(_0507_),
    .Y(_1196_)
  );
  NAND _1278_ (
    .A(_1170_),
    .B(_1175_),
    .Y(_0508_)
  );
  NOR _1279_ (
    .A(_0463_),
    .B(_0479_),
    .Y(_0509_)
  );
  NOR _1280_ (
    .A(_0971_),
    .B(_0982_),
    .Y(_0510_)
  );
  NAND _1281_ (
    .A(_0463_),
    .B(_0479_),
    .Y(_0511_)
  );
  NOR _1282_ (
    .A(_0509_),
    .B(_0510_),
    .Y(_0512_)
  );
  NOR _1283_ (
    .A(_0508_),
    .B(_0512_),
    .Y(_0513_)
  );
  NAND _1284_ (
    .A(_0508_),
    .B(_0512_),
    .Y(_0514_)
  );
  NAND _1285_ (
    .A(_1178_),
    .B(_0514_),
    .Y(_0515_)
  );
  NOR _1286_ (
    .A(_0513_),
    .B(_0515_),
    .Y(_0516_)
  );
  NOR _1287_ (
    .A(_0463_),
    .B(_0480_),
    .Y(_0517_)
  );
  NAND _1288_ (
    .A(_0463_),
    .B(_0480_),
    .Y(_0518_)
  );
  NOT _1289_ (
    .A(_0518_),
    .Y(_0519_)
  );
  NOR _1290_ (
    .A(_0517_),
    .B(_0519_),
    .Y(_0520_)
  );
  NOR _1291_ (
    .A(_0500_),
    .B(_0520_),
    .Y(_0521_)
  );
  NAND _1292_ (
    .A(_0500_),
    .B(_0520_),
    .Y(_0522_)
  );
  NAND _1293_ (
    .A(_0498_),
    .B(_0522_),
    .Y(_0523_)
  );
  NOR _1294_ (
    .A(_0521_),
    .B(_0523_),
    .Y(_0524_)
  );
  NAND _1295_ (
    .A(_0463_),
    .B(_0464_),
    .Y(_0525_)
  );
  NOR _1296_ (
    .A(_0456_),
    .B(_0525_),
    .Y(_0526_)
  );
  NOR _1297_ (
    .A(_0456_),
    .B(_0971_),
    .Y(_0527_)
  );
  NOR _1298_ (
    .A(_0464_),
    .B(_0527_),
    .Y(_0528_)
  );
  NOR _1299_ (
    .A(_0492_),
    .B(_0528_),
    .Y(_0529_)
  );
  NOT _1300_ (
    .A(_0529_),
    .Y(_0530_)
  );
  NOR _1301_ (
    .A(_0526_),
    .B(_0530_),
    .Y(_0531_)
  );
  NOR _1302_ (
    .A(_1191_),
    .B(_0509_),
    .Y(_0532_)
  );
  NOR _1303_ (
    .A(_1183_),
    .B(_0511_),
    .Y(_0533_)
  );
  NOT _1304_ (
    .A(_0533_),
    .Y(_0534_)
  );
  NAND _1305_ (
    .A(_1195_),
    .B(_1185_),
    .Y(_0535_)
  );
  NOR _1306_ (
    .A(_0463_),
    .B(_0535_),
    .Y(_0536_)
  );
  NOT _1307_ (
    .A(_0536_),
    .Y(_0537_)
  );
  NOR _1308_ (
    .A(_1195_),
    .B(_1186_),
    .Y(_0538_)
  );
  NAND _1309_ (
    .A(_0950_),
    .B(_1185_),
    .Y(_0539_)
  );
  NAND _1310_ (
    .A(_0496_),
    .B(_0538_),
    .Y(_0540_)
  );
  NOR _1311_ (
    .A(_0516_),
    .B(_0532_),
    .Y(_0541_)
  );
  NOR _1312_ (
    .A(_0524_),
    .B(_0531_),
    .Y(_0542_)
  );
  NAND _1313_ (
    .A(_0537_),
    .B(_0542_),
    .Y(_0543_)
  );
  NAND _1314_ (
    .A(_0534_),
    .B(_0540_),
    .Y(_0544_)
  );
  NOR _1315_ (
    .A(_0543_),
    .B(_0544_),
    .Y(_0545_)
  );
  NAND _1316_ (
    .A(_0541_),
    .B(_0545_),
    .Y(_1202_)
  );
  NOT _1317_ (
    .A(_1202_),
    .Y(_0546_)
  );
  NAND _1318_ (
    .A(_0511_),
    .B(_0514_),
    .Y(_0547_)
  );
  NOR _1319_ (
    .A(_0993_),
    .B(_1004_),
    .Y(_0548_)
  );
  NAND _1320_ (
    .A(_0464_),
    .B(_0480_),
    .Y(_0549_)
  );
  NOR _1321_ (
    .A(_0464_),
    .B(_0480_),
    .Y(_0550_)
  );
  NOR _1322_ (
    .A(_0548_),
    .B(_0550_),
    .Y(_0551_)
  );
  NOR _1323_ (
    .A(_0547_),
    .B(_0551_),
    .Y(_0552_)
  );
  NAND _1324_ (
    .A(_0547_),
    .B(_0551_),
    .Y(_0553_)
  );
  NOR _1325_ (
    .A(_1179_),
    .B(_0552_),
    .Y(_0554_)
  );
  NAND _1326_ (
    .A(_0553_),
    .B(_0554_),
    .Y(_0555_)
  );
  NAND _1327_ (
    .A(_0518_),
    .B(_0522_),
    .Y(_0556_)
  );
  NOT _1328_ (
    .A(_0556_),
    .Y(_0557_)
  );
  NAND _1329_ (
    .A(_0464_),
    .B(_0481_),
    .Y(_0558_)
  );
  NOR _1330_ (
    .A(_0464_),
    .B(_0481_),
    .Y(_0559_)
  );
  NOT _1331_ (
    .A(_0559_),
    .Y(_0560_)
  );
  NAND _1332_ (
    .A(_0558_),
    .B(_0560_),
    .Y(_0561_)
  );
  NOT _1333_ (
    .A(_0561_),
    .Y(_0562_)
  );
  NAND _1334_ (
    .A(_0556_),
    .B(_0562_),
    .Y(_0563_)
  );
  NAND _1335_ (
    .A(_0557_),
    .B(_0561_),
    .Y(_0564_)
  );
  NAND _1336_ (
    .A(_0563_),
    .B(_0564_),
    .Y(_0565_)
  );
  NOR _1337_ (
    .A(_0499_),
    .B(_0565_),
    .Y(_0566_)
  );
  NOR _1338_ (
    .A(_0464_),
    .B(_0465_),
    .Y(_0567_)
  );
  NAND _1339_ (
    .A(_0464_),
    .B(_0465_),
    .Y(_0568_)
  );
  NOT _1340_ (
    .A(_0568_),
    .Y(_0569_)
  );
  NOR _1341_ (
    .A(_0567_),
    .B(_0569_),
    .Y(_0570_)
  );
  NAND _1342_ (
    .A(_0494_),
    .B(_0525_),
    .Y(_0571_)
  );
  NOR _1343_ (
    .A(_0570_),
    .B(_0571_),
    .Y(_0572_)
  );
  NAND _1344_ (
    .A(_0570_),
    .B(_0571_),
    .Y(_0573_)
  );
  NAND _1345_ (
    .A(_0491_),
    .B(_0573_),
    .Y(_0574_)
  );
  NOR _1346_ (
    .A(_0572_),
    .B(_0574_),
    .Y(_0575_)
  );
  NAND _1347_ (
    .A(_0993_),
    .B(_0494_),
    .Y(_0576_)
  );
  NOR _1348_ (
    .A(_0993_),
    .B(_0494_),
    .Y(_0577_)
  );
  NOR _1349_ (
    .A(_0539_),
    .B(_0577_),
    .Y(_0578_)
  );
  NAND _1350_ (
    .A(_0576_),
    .B(_0578_),
    .Y(_0579_)
  );
  NOR _1351_ (
    .A(_1191_),
    .B(_0550_),
    .Y(_0580_)
  );
  NOR _1352_ (
    .A(_0464_),
    .B(_0535_),
    .Y(_0581_)
  );
  NOR _1353_ (
    .A(_1183_),
    .B(_0549_),
    .Y(_0582_)
  );
  NOT _1354_ (
    .A(_0582_),
    .Y(_0583_)
  );
  NOR _1355_ (
    .A(_0580_),
    .B(_0581_),
    .Y(_0584_)
  );
  NAND _1356_ (
    .A(_0579_),
    .B(_0584_),
    .Y(_0585_)
  );
  NOR _1357_ (
    .A(_0575_),
    .B(_0585_),
    .Y(_0586_)
  );
  NAND _1358_ (
    .A(_0583_),
    .B(_0586_),
    .Y(_0587_)
  );
  NOR _1359_ (
    .A(_0566_),
    .B(_0587_),
    .Y(_0588_)
  );
  NAND _1360_ (
    .A(_0555_),
    .B(_0588_),
    .Y(_1203_)
  );
  NAND _1361_ (
    .A(_0549_),
    .B(_0553_),
    .Y(_0589_)
  );
  NOR _1362_ (
    .A(_0465_),
    .B(_0481_),
    .Y(_0590_)
  );
  NOR _1363_ (
    .A(_1015_),
    .B(_1025_),
    .Y(_0591_)
  );
  NAND _1364_ (
    .A(_0465_),
    .B(_0481_),
    .Y(_0592_)
  );
  NOR _1365_ (
    .A(_0590_),
    .B(_0591_),
    .Y(_0593_)
  );
  NOR _1366_ (
    .A(_0589_),
    .B(_0593_),
    .Y(_0594_)
  );
  NAND _1367_ (
    .A(_0589_),
    .B(_0593_),
    .Y(_0595_)
  );
  NOR _1368_ (
    .A(_1179_),
    .B(_0594_),
    .Y(_0596_)
  );
  NAND _1369_ (
    .A(_0595_),
    .B(_0596_),
    .Y(_0597_)
  );
  NAND _1370_ (
    .A(_0558_),
    .B(_0563_),
    .Y(_0598_)
  );
  NOR _1371_ (
    .A(_0465_),
    .B(_0482_),
    .Y(_0599_)
  );
  NOR _1372_ (
    .A(_1015_),
    .B(_1036_),
    .Y(_0600_)
  );
  NOR _1373_ (
    .A(_0599_),
    .B(_0600_),
    .Y(_0601_)
  );
  NAND _1374_ (
    .A(_0598_),
    .B(_0601_),
    .Y(_0602_)
  );
  NOR _1375_ (
    .A(_0598_),
    .B(_0601_),
    .Y(_0603_)
  );
  NAND _1376_ (
    .A(_0498_),
    .B(_0602_),
    .Y(_0604_)
  );
  NOR _1377_ (
    .A(_0603_),
    .B(_0604_),
    .Y(_0605_)
  );
  NAND _1378_ (
    .A(_0568_),
    .B(_0573_),
    .Y(_0606_)
  );
  NOR _1379_ (
    .A(_0465_),
    .B(_0466_),
    .Y(_0607_)
  );
  NOT _1380_ (
    .A(_0607_),
    .Y(_0608_)
  );
  NAND _1381_ (
    .A(_0465_),
    .B(_0466_),
    .Y(_0609_)
  );
  NOT _1382_ (
    .A(_0609_),
    .Y(_0610_)
  );
  NOR _1383_ (
    .A(_0607_),
    .B(_0610_),
    .Y(_0611_)
  );
  NAND _1384_ (
    .A(_0606_),
    .B(_0611_),
    .Y(_0612_)
  );
  NOR _1385_ (
    .A(_0606_),
    .B(_0611_),
    .Y(_0613_)
  );
  NOR _1386_ (
    .A(_0492_),
    .B(_0613_),
    .Y(_0614_)
  );
  NAND _1387_ (
    .A(_0612_),
    .B(_0614_),
    .Y(_0615_)
  );
  NOR _1388_ (
    .A(_0465_),
    .B(_0577_),
    .Y(_0616_)
  );
  NOR _1389_ (
    .A(_0494_),
    .B(_0568_),
    .Y(_0617_)
  );
  NOR _1390_ (
    .A(_0616_),
    .B(_0617_),
    .Y(_0618_)
  );
  NAND _1391_ (
    .A(_0538_),
    .B(_0618_),
    .Y(_0619_)
  );
  NOR _1392_ (
    .A(_0465_),
    .B(_0535_),
    .Y(_0620_)
  );
  NOR _1393_ (
    .A(_1191_),
    .B(_0590_),
    .Y(_0621_)
  );
  NOR _1394_ (
    .A(_1183_),
    .B(_0592_),
    .Y(_0622_)
  );
  NOR _1395_ (
    .A(_0620_),
    .B(_0622_),
    .Y(_0623_)
  );
  NAND _1396_ (
    .A(_0619_),
    .B(_0623_),
    .Y(_0624_)
  );
  NOR _1397_ (
    .A(_0621_),
    .B(_0624_),
    .Y(_0625_)
  );
  NAND _1398_ (
    .A(_0615_),
    .B(_0625_),
    .Y(_0626_)
  );
  NOR _1399_ (
    .A(_0605_),
    .B(_0626_),
    .Y(_0627_)
  );
  NAND _1400_ (
    .A(_0597_),
    .B(_0627_),
    .Y(_1204_)
  );
  NAND _1401_ (
    .A(_0466_),
    .B(_0482_),
    .Y(_0628_)
  );
  NOT _1402_ (
    .A(_0628_),
    .Y(_0629_)
  );
  NOR _1403_ (
    .A(_0466_),
    .B(_0482_),
    .Y(_0630_)
  );
  NOR _1404_ (
    .A(_0629_),
    .B(_0630_),
    .Y(_0631_)
  );
  NOR _1405_ (
    .A(_0589_),
    .B(_0591_),
    .Y(_0632_)
  );
  NOR _1406_ (
    .A(_0590_),
    .B(_0632_),
    .Y(_0633_)
  );
  NOR _1407_ (
    .A(_0631_),
    .B(_0633_),
    .Y(_0634_)
  );
  NAND _1408_ (
    .A(_0631_),
    .B(_0633_),
    .Y(_0635_)
  );
  NOR _1409_ (
    .A(_1179_),
    .B(_0634_),
    .Y(_0636_)
  );
  NAND _1410_ (
    .A(_0635_),
    .B(_0636_),
    .Y(_0637_)
  );
  NAND _1411_ (
    .A(_0466_),
    .B(_0483_),
    .Y(_0638_)
  );
  NOT _1412_ (
    .A(_0638_),
    .Y(_0639_)
  );
  NOR _1413_ (
    .A(_0466_),
    .B(_0483_),
    .Y(_0640_)
  );
  NOR _1414_ (
    .A(_0639_),
    .B(_0640_),
    .Y(_0641_)
  );
  NOR _1415_ (
    .A(_0598_),
    .B(_0600_),
    .Y(_0642_)
  );
  NOR _1416_ (
    .A(_0599_),
    .B(_0642_),
    .Y(_0643_)
  );
  NOR _1417_ (
    .A(_0641_),
    .B(_0643_),
    .Y(_0644_)
  );
  NAND _1418_ (
    .A(_0641_),
    .B(_0643_),
    .Y(_0645_)
  );
  NAND _1419_ (
    .A(_0498_),
    .B(_0645_),
    .Y(_0646_)
  );
  NOR _1420_ (
    .A(_0644_),
    .B(_0646_),
    .Y(_0647_)
  );
  NOR _1421_ (
    .A(_0466_),
    .B(_0617_),
    .Y(_0648_)
  );
  NAND _1422_ (
    .A(_0466_),
    .B(_0617_),
    .Y(_0649_)
  );
  NOT _1423_ (
    .A(_0649_),
    .Y(_0650_)
  );
  NAND _1424_ (
    .A(_0538_),
    .B(_0649_),
    .Y(_0651_)
  );
  NOR _1425_ (
    .A(_0648_),
    .B(_0651_),
    .Y(_0652_)
  );
  NOT _1426_ (
    .A(_0652_),
    .Y(_0653_)
  );
  NOR _1427_ (
    .A(_1191_),
    .B(_0630_),
    .Y(_0654_)
  );
  NOR _1428_ (
    .A(_1183_),
    .B(_0628_),
    .Y(_0655_)
  );
  NOR _1429_ (
    .A(_0466_),
    .B(_0535_),
    .Y(_0656_)
  );
  NOR _1430_ (
    .A(_0654_),
    .B(_0656_),
    .Y(_0657_)
  );
  NAND _1431_ (
    .A(_0653_),
    .B(_0657_),
    .Y(_0658_)
  );
  NOR _1432_ (
    .A(_0655_),
    .B(_0658_),
    .Y(_0659_)
  );
  NAND _1433_ (
    .A(_0573_),
    .B(_0609_),
    .Y(_0660_)
  );
  NAND _1434_ (
    .A(_0608_),
    .B(_0660_),
    .Y(_0661_)
  );
  NAND _1435_ (
    .A(_0568_),
    .B(_0661_),
    .Y(_0662_)
  );
  NOR _1436_ (
    .A(_0466_),
    .B(_0467_),
    .Y(_0663_)
  );
  NAND _1437_ (
    .A(_0466_),
    .B(_0467_),
    .Y(_0664_)
  );
  NOT _1438_ (
    .A(_0664_),
    .Y(_0665_)
  );
  NOR _1439_ (
    .A(_0663_),
    .B(_0665_),
    .Y(_0666_)
  );
  NAND _1440_ (
    .A(_0662_),
    .B(_0666_),
    .Y(_0667_)
  );
  NOR _1441_ (
    .A(_0662_),
    .B(_0666_),
    .Y(_0668_)
  );
  NOR _1442_ (
    .A(_0492_),
    .B(_0668_),
    .Y(_0669_)
  );
  NAND _1443_ (
    .A(_0667_),
    .B(_0669_),
    .Y(_0670_)
  );
  NAND _1444_ (
    .A(_0659_),
    .B(_0670_),
    .Y(_0671_)
  );
  NOR _1445_ (
    .A(_0647_),
    .B(_0671_),
    .Y(_0672_)
  );
  NAND _1446_ (
    .A(_0637_),
    .B(_0672_),
    .Y(_1205_)
  );
  NAND _1447_ (
    .A(_0628_),
    .B(_0635_),
    .Y(_0673_)
  );
  NAND _1448_ (
    .A(_0467_),
    .B(_0483_),
    .Y(_0674_)
  );
  NOT _1449_ (
    .A(_0674_),
    .Y(_0675_)
  );
  NOR _1450_ (
    .A(_0467_),
    .B(_0483_),
    .Y(_0676_)
  );
  NOR _1451_ (
    .A(_0675_),
    .B(_0676_),
    .Y(_0677_)
  );
  NAND _1452_ (
    .A(_0673_),
    .B(_0677_),
    .Y(_0678_)
  );
  NOR _1453_ (
    .A(_0673_),
    .B(_0677_),
    .Y(_0679_)
  );
  NOR _1454_ (
    .A(_1179_),
    .B(_0679_),
    .Y(_0680_)
  );
  NAND _1455_ (
    .A(_0678_),
    .B(_0680_),
    .Y(_0681_)
  );
  NAND _1456_ (
    .A(_0638_),
    .B(_0645_),
    .Y(_0682_)
  );
  NOR _1457_ (
    .A(_0467_),
    .B(_0484_),
    .Y(_0683_)
  );
  NAND _1458_ (
    .A(_0467_),
    .B(_0484_),
    .Y(_0684_)
  );
  NOT _1459_ (
    .A(_0684_),
    .Y(_0685_)
  );
  NOR _1460_ (
    .A(_0683_),
    .B(_0685_),
    .Y(_0686_)
  );
  NAND _1461_ (
    .A(_0682_),
    .B(_0686_),
    .Y(_0687_)
  );
  NOR _1462_ (
    .A(_0682_),
    .B(_0686_),
    .Y(_0688_)
  );
  NAND _1463_ (
    .A(_0498_),
    .B(_0687_),
    .Y(_0689_)
  );
  NOR _1464_ (
    .A(_0688_),
    .B(_0689_),
    .Y(_0690_)
  );
  NAND _1465_ (
    .A(_0664_),
    .B(_0667_),
    .Y(_0691_)
  );
  NOR _1466_ (
    .A(_0467_),
    .B(_0468_),
    .Y(_0692_)
  );
  NOT _1467_ (
    .A(_0692_),
    .Y(_0693_)
  );
  NAND _1468_ (
    .A(_0467_),
    .B(_0468_),
    .Y(_0694_)
  );
  NOT _1469_ (
    .A(_0694_),
    .Y(_0695_)
  );
  NOR _1470_ (
    .A(_0692_),
    .B(_0695_),
    .Y(_0696_)
  );
  NOR _1471_ (
    .A(_0691_),
    .B(_0696_),
    .Y(_0697_)
  );
  NAND _1472_ (
    .A(_0691_),
    .B(_0696_),
    .Y(_0698_)
  );
  NOR _1473_ (
    .A(_0492_),
    .B(_0697_),
    .Y(_0699_)
  );
  NAND _1474_ (
    .A(_0698_),
    .B(_0699_),
    .Y(_0700_)
  );
  NOR _1475_ (
    .A(_0467_),
    .B(_0650_),
    .Y(_0701_)
  );
  NAND _1476_ (
    .A(_0467_),
    .B(_0650_),
    .Y(_0702_)
  );
  NAND _1477_ (
    .A(_0538_),
    .B(_0702_),
    .Y(_0703_)
  );
  NOR _1478_ (
    .A(_0701_),
    .B(_0703_),
    .Y(_0704_)
  );
  NOR _1479_ (
    .A(_1191_),
    .B(_0676_),
    .Y(_0705_)
  );
  NOR _1480_ (
    .A(_0467_),
    .B(_0535_),
    .Y(_0706_)
  );
  NAND _1481_ (
    .A(_1182_),
    .B(_0675_),
    .Y(_0707_)
  );
  NOR _1482_ (
    .A(_0705_),
    .B(_0706_),
    .Y(_0708_)
  );
  NAND _1483_ (
    .A(_0707_),
    .B(_0708_),
    .Y(_0709_)
  );
  NOR _1484_ (
    .A(_0704_),
    .B(_0709_),
    .Y(_0710_)
  );
  NAND _1485_ (
    .A(_0700_),
    .B(_0710_),
    .Y(_0711_)
  );
  NOR _1486_ (
    .A(_0690_),
    .B(_0711_),
    .Y(_0712_)
  );
  NAND _1487_ (
    .A(_0681_),
    .B(_0712_),
    .Y(_1206_)
  );
  NAND _1488_ (
    .A(_0674_),
    .B(_0678_),
    .Y(_0713_)
  );
  NAND _1489_ (
    .A(_0468_),
    .B(_0484_),
    .Y(_0714_)
  );
  NOT _1490_ (
    .A(_0714_),
    .Y(_0715_)
  );
  NOR _1491_ (
    .A(_0468_),
    .B(_0484_),
    .Y(_0716_)
  );
  NOR _1492_ (
    .A(_0715_),
    .B(_0716_),
    .Y(_0717_)
  );
  NAND _1493_ (
    .A(_0713_),
    .B(_0717_),
    .Y(_0718_)
  );
  NOR _1494_ (
    .A(_0713_),
    .B(_0717_),
    .Y(_0719_)
  );
  NOR _1495_ (
    .A(_1179_),
    .B(_0719_),
    .Y(_0720_)
  );
  NAND _1496_ (
    .A(_0718_),
    .B(_0720_),
    .Y(_0721_)
  );
  NAND _1497_ (
    .A(_0684_),
    .B(_0687_),
    .Y(_0722_)
  );
  NOR _1498_ (
    .A(_0468_),
    .B(_0485_),
    .Y(_0723_)
  );
  NAND _1499_ (
    .A(_0468_),
    .B(_0485_),
    .Y(_0724_)
  );
  NOT _1500_ (
    .A(_0724_),
    .Y(_0725_)
  );
  NOR _1501_ (
    .A(_0723_),
    .B(_0725_),
    .Y(_0726_)
  );
  NOR _1502_ (
    .A(_0722_),
    .B(_0726_),
    .Y(_0727_)
  );
  NAND _1503_ (
    .A(_0722_),
    .B(_0726_),
    .Y(_0728_)
  );
  NAND _1504_ (
    .A(_0498_),
    .B(_0728_),
    .Y(_0729_)
  );
  NOR _1505_ (
    .A(_0727_),
    .B(_0729_),
    .Y(_0730_)
  );
  NAND _1506_ (
    .A(_0667_),
    .B(_0694_),
    .Y(_0731_)
  );
  NAND _1507_ (
    .A(_0693_),
    .B(_0731_),
    .Y(_0732_)
  );
  NAND _1508_ (
    .A(_0664_),
    .B(_0732_),
    .Y(_0733_)
  );
  NAND _1509_ (
    .A(_0468_),
    .B(_0469_),
    .Y(_0734_)
  );
  NOT _1510_ (
    .A(_0734_),
    .Y(_0735_)
  );
  NOR _1511_ (
    .A(_0468_),
    .B(_0469_),
    .Y(_0736_)
  );
  NOR _1512_ (
    .A(_0735_),
    .B(_0736_),
    .Y(_0737_)
  );
  NOR _1513_ (
    .A(_0733_),
    .B(_0737_),
    .Y(_0738_)
  );
  NAND _1514_ (
    .A(_0733_),
    .B(_0737_),
    .Y(_0739_)
  );
  NOT _1515_ (
    .A(_0739_),
    .Y(_0740_)
  );
  NOR _1516_ (
    .A(_0738_),
    .B(_0740_),
    .Y(_0741_)
  );
  NAND _1517_ (
    .A(_0491_),
    .B(_0741_),
    .Y(_0742_)
  );
  NAND _1518_ (
    .A(_1047_),
    .B(_0702_),
    .Y(_0743_)
  );
  NOR _1519_ (
    .A(_0649_),
    .B(_0694_),
    .Y(_0744_)
  );
  NOR _1520_ (
    .A(_0539_),
    .B(_0744_),
    .Y(_0745_)
  );
  NAND _1521_ (
    .A(_0743_),
    .B(_0745_),
    .Y(_0746_)
  );
  NOR _1522_ (
    .A(_1191_),
    .B(_0716_),
    .Y(_0747_)
  );
  NOR _1523_ (
    .A(_1183_),
    .B(_0714_),
    .Y(_0748_)
  );
  NOR _1524_ (
    .A(_0468_),
    .B(_0535_),
    .Y(_0749_)
  );
  NOR _1525_ (
    .A(_0747_),
    .B(_0749_),
    .Y(_0750_)
  );
  NAND _1526_ (
    .A(_0746_),
    .B(_0750_),
    .Y(_0751_)
  );
  NOR _1527_ (
    .A(_0748_),
    .B(_0751_),
    .Y(_0752_)
  );
  NAND _1528_ (
    .A(_0742_),
    .B(_0752_),
    .Y(_0753_)
  );
  NOR _1529_ (
    .A(_0730_),
    .B(_0753_),
    .Y(_0754_)
  );
  NAND _1530_ (
    .A(_0721_),
    .B(_0754_),
    .Y(_1207_)
  );
  NAND _1531_ (
    .A(_0714_),
    .B(_0718_),
    .Y(_0755_)
  );
  NAND _1532_ (
    .A(_0469_),
    .B(_0485_),
    .Y(_0756_)
  );
  NOT _1533_ (
    .A(_0756_),
    .Y(_0757_)
  );
  NOR _1534_ (
    .A(_0469_),
    .B(_0485_),
    .Y(_0758_)
  );
  NOR _1535_ (
    .A(_0757_),
    .B(_0758_),
    .Y(_0759_)
  );
  NAND _1536_ (
    .A(_0755_),
    .B(_0759_),
    .Y(_0760_)
  );
  NOR _1537_ (
    .A(_0755_),
    .B(_0759_),
    .Y(_0761_)
  );
  NOR _1538_ (
    .A(_1179_),
    .B(_0761_),
    .Y(_0762_)
  );
  NAND _1539_ (
    .A(_0760_),
    .B(_0762_),
    .Y(_0763_)
  );
  NAND _1540_ (
    .A(_0724_),
    .B(_0728_),
    .Y(_0764_)
  );
  NOR _1541_ (
    .A(_0469_),
    .B(_0486_),
    .Y(_0765_)
  );
  NOR _1542_ (
    .A(_1058_),
    .B(_1079_),
    .Y(_0766_)
  );
  NOR _1543_ (
    .A(_0765_),
    .B(_0766_),
    .Y(_0767_)
  );
  NOR _1544_ (
    .A(_0764_),
    .B(_0767_),
    .Y(_0768_)
  );
  NAND _1545_ (
    .A(_0764_),
    .B(_0767_),
    .Y(_0769_)
  );
  NOR _1546_ (
    .A(_0499_),
    .B(_0768_),
    .Y(_0770_)
  );
  NAND _1547_ (
    .A(_0769_),
    .B(_0770_),
    .Y(_0771_)
  );
  NOR _1548_ (
    .A(_0469_),
    .B(_0744_),
    .Y(_0772_)
  );
  NOR _1549_ (
    .A(_0702_),
    .B(_0734_),
    .Y(_0773_)
  );
  NAND _1550_ (
    .A(_0469_),
    .B(_0744_),
    .Y(_0774_)
  );
  NOT _1551_ (
    .A(_0774_),
    .Y(_0775_)
  );
  NOR _1552_ (
    .A(_0772_),
    .B(_0775_),
    .Y(_0776_)
  );
  NAND _1553_ (
    .A(_0538_),
    .B(_0776_),
    .Y(_0777_)
  );
  NOR _1554_ (
    .A(_1191_),
    .B(_0758_),
    .Y(_0778_)
  );
  NOR _1555_ (
    .A(_1183_),
    .B(_0756_),
    .Y(_0779_)
  );
  NOR _1556_ (
    .A(_0469_),
    .B(_0535_),
    .Y(_0780_)
  );
  NOR _1557_ (
    .A(_0778_),
    .B(_0779_),
    .Y(_0781_)
  );
  NOT _1558_ (
    .A(_0781_),
    .Y(_0782_)
  );
  NOR _1559_ (
    .A(_0780_),
    .B(_0782_),
    .Y(_0783_)
  );
  NAND _1560_ (
    .A(_0777_),
    .B(_0783_),
    .Y(_0784_)
  );
  NAND _1561_ (
    .A(_0734_),
    .B(_0739_),
    .Y(_0785_)
  );
  NOR _1562_ (
    .A(_0469_),
    .B(_0470_),
    .Y(_0786_)
  );
  NAND _1563_ (
    .A(_0469_),
    .B(_0470_),
    .Y(_0787_)
  );
  NOT _1564_ (
    .A(_0787_),
    .Y(_0788_)
  );
  NOR _1565_ (
    .A(_0786_),
    .B(_0788_),
    .Y(_0789_)
  );
  NAND _1566_ (
    .A(_0785_),
    .B(_0789_),
    .Y(_0790_)
  );
  NOR _1567_ (
    .A(_0785_),
    .B(_0789_),
    .Y(_0791_)
  );
  NOR _1568_ (
    .A(_0492_),
    .B(_0791_),
    .Y(_0792_)
  );
  NAND _1569_ (
    .A(_0790_),
    .B(_0792_),
    .Y(_0793_)
  );
  NAND _1570_ (
    .A(_0771_),
    .B(_0793_),
    .Y(_0794_)
  );
  NOR _1571_ (
    .A(_0784_),
    .B(_0794_),
    .Y(_0795_)
  );
  NAND _1572_ (
    .A(_0763_),
    .B(_0795_),
    .Y(_1208_)
  );
  NOR _1573_ (
    .A(_1069_),
    .B(_1079_),
    .Y(_0796_)
  );
  NAND _1574_ (
    .A(_0470_),
    .B(_0486_),
    .Y(_0797_)
  );
  NOR _1575_ (
    .A(_0470_),
    .B(_0486_),
    .Y(_0798_)
  );
  NOR _1576_ (
    .A(_0796_),
    .B(_0798_),
    .Y(_0799_)
  );
  NOR _1577_ (
    .A(_0755_),
    .B(_0757_),
    .Y(_0800_)
  );
  NOR _1578_ (
    .A(_0758_),
    .B(_0800_),
    .Y(_0801_)
  );
  NAND _1579_ (
    .A(_0799_),
    .B(_0801_),
    .Y(_0802_)
  );
  NOR _1580_ (
    .A(_0799_),
    .B(_0801_),
    .Y(_0803_)
  );
  NOR _1581_ (
    .A(_1179_),
    .B(_0803_),
    .Y(_0804_)
  );
  NAND _1582_ (
    .A(_0802_),
    .B(_0804_),
    .Y(_0805_)
  );
  NOR _1583_ (
    .A(_0470_),
    .B(_0487_),
    .Y(_0806_)
  );
  NAND _1584_ (
    .A(_0470_),
    .B(_0487_),
    .Y(_0807_)
  );
  NOT _1585_ (
    .A(_0807_),
    .Y(_0808_)
  );
  NOR _1586_ (
    .A(_0806_),
    .B(_0808_),
    .Y(_0809_)
  );
  NOR _1587_ (
    .A(_0764_),
    .B(_0766_),
    .Y(_0810_)
  );
  NOR _1588_ (
    .A(_0765_),
    .B(_0810_),
    .Y(_0811_)
  );
  NOR _1589_ (
    .A(_0809_),
    .B(_0811_),
    .Y(_0812_)
  );
  NAND _1590_ (
    .A(_0809_),
    .B(_0811_),
    .Y(_0813_)
  );
  NAND _1591_ (
    .A(_0498_),
    .B(_0813_),
    .Y(_0814_)
  );
  NOR _1592_ (
    .A(_0812_),
    .B(_0814_),
    .Y(_0815_)
  );
  NOR _1593_ (
    .A(_0470_),
    .B(_0775_),
    .Y(_0816_)
  );
  NAND _1594_ (
    .A(_0744_),
    .B(_0788_),
    .Y(_0817_)
  );
  NOT _1595_ (
    .A(_0817_),
    .Y(_0818_)
  );
  NAND _1596_ (
    .A(_0538_),
    .B(_0817_),
    .Y(_0819_)
  );
  NOR _1597_ (
    .A(_0816_),
    .B(_0819_),
    .Y(_0820_)
  );
  NOR _1598_ (
    .A(_1191_),
    .B(_0798_),
    .Y(_0821_)
  );
  NAND _1599_ (
    .A(_1182_),
    .B(_0796_),
    .Y(_0822_)
  );
  NOR _1600_ (
    .A(_0470_),
    .B(_0535_),
    .Y(_0823_)
  );
  NOR _1601_ (
    .A(_0821_),
    .B(_0823_),
    .Y(_0824_)
  );
  NAND _1602_ (
    .A(_0822_),
    .B(_0824_),
    .Y(_0825_)
  );
  NOR _1603_ (
    .A(_0820_),
    .B(_0825_),
    .Y(_0826_)
  );
  NAND _1604_ (
    .A(_0740_),
    .B(_0789_),
    .Y(_0827_)
  );
  NAND _1605_ (
    .A(_0787_),
    .B(_0827_),
    .Y(_0828_)
  );
  NOR _1606_ (
    .A(_0735_),
    .B(_0828_),
    .Y(_0829_)
  );
  NAND _1607_ (
    .A(_0470_),
    .B(_0471_),
    .Y(_0830_)
  );
  NOT _1608_ (
    .A(_0830_),
    .Y(_0831_)
  );
  NOR _1609_ (
    .A(_0470_),
    .B(_0471_),
    .Y(_0832_)
  );
  NOT _1610_ (
    .A(_0832_),
    .Y(_0833_)
  );
  NAND _1611_ (
    .A(_0830_),
    .B(_0833_),
    .Y(_0834_)
  );
  NAND _1612_ (
    .A(_0829_),
    .B(_0834_),
    .Y(_0835_)
  );
  NOR _1613_ (
    .A(_0829_),
    .B(_0834_),
    .Y(_0836_)
  );
  NOT _1614_ (
    .A(_0836_),
    .Y(_0837_)
  );
  NOR _1615_ (
    .A(_0492_),
    .B(_0836_),
    .Y(_0838_)
  );
  NAND _1616_ (
    .A(_0835_),
    .B(_0838_),
    .Y(_0839_)
  );
  NAND _1617_ (
    .A(_0826_),
    .B(_0839_),
    .Y(_0840_)
  );
  NOR _1618_ (
    .A(_0815_),
    .B(_0840_),
    .Y(_0841_)
  );
  NAND _1619_ (
    .A(_0805_),
    .B(_0841_),
    .Y(_1209_)
  );
  NAND _1620_ (
    .A(_0797_),
    .B(_0802_),
    .Y(_0842_)
  );
  NOR _1621_ (
    .A(_0471_),
    .B(_0487_),
    .Y(_0843_)
  );
  NAND _1622_ (
    .A(_0471_),
    .B(_0487_),
    .Y(_0844_)
  );
  NOT _1623_ (
    .A(_0844_),
    .Y(_0845_)
  );
  NOR _1624_ (
    .A(_0843_),
    .B(_0845_),
    .Y(_0846_)
  );
  NAND _1625_ (
    .A(_0842_),
    .B(_0846_),
    .Y(_0847_)
  );
  NOR _1626_ (
    .A(_0842_),
    .B(_0846_),
    .Y(_0848_)
  );
  NOR _1627_ (
    .A(_1179_),
    .B(_0848_),
    .Y(_0849_)
  );
  NAND _1628_ (
    .A(_0847_),
    .B(_0849_),
    .Y(_0850_)
  );
  NAND _1629_ (
    .A(_0807_),
    .B(_0813_),
    .Y(_0851_)
  );
  NOT _1630_ (
    .A(_0851_),
    .Y(_0852_)
  );
  NAND _1631_ (
    .A(_1090_),
    .B(_1112_),
    .Y(_0853_)
  );
  NAND _1632_ (
    .A(_0471_),
    .B(_0473_),
    .Y(_0854_)
  );
  NAND _1633_ (
    .A(_0853_),
    .B(_0854_),
    .Y(_0855_)
  );
  NOR _1634_ (
    .A(_0852_),
    .B(_0855_),
    .Y(_0856_)
  );
  NAND _1635_ (
    .A(_0852_),
    .B(_0855_),
    .Y(_0857_)
  );
  NAND _1636_ (
    .A(_0498_),
    .B(_0857_),
    .Y(_0858_)
  );
  NOR _1637_ (
    .A(_0856_),
    .B(_0858_),
    .Y(_0859_)
  );
  NAND _1638_ (
    .A(_1090_),
    .B(_0817_),
    .Y(_0860_)
  );
  NAND _1639_ (
    .A(_0773_),
    .B(_0831_),
    .Y(_0861_)
  );
  NOR _1640_ (
    .A(_0774_),
    .B(_0830_),
    .Y(_0862_)
  );
  NOR _1641_ (
    .A(_0539_),
    .B(_0862_),
    .Y(_0863_)
  );
  NAND _1642_ (
    .A(_0860_),
    .B(_0863_),
    .Y(_0864_)
  );
  NOR _1643_ (
    .A(_0471_),
    .B(_0535_),
    .Y(_0865_)
  );
  NOR _1644_ (
    .A(_1183_),
    .B(_0844_),
    .Y(_0866_)
  );
  NOR _1645_ (
    .A(_1191_),
    .B(_0843_),
    .Y(_0867_)
  );
  NOR _1646_ (
    .A(_0865_),
    .B(_0867_),
    .Y(_0868_)
  );
  NAND _1647_ (
    .A(_0864_),
    .B(_0868_),
    .Y(_0869_)
  );
  NOR _1648_ (
    .A(_0866_),
    .B(_0869_),
    .Y(_0870_)
  );
  NAND _1649_ (
    .A(_0830_),
    .B(_0837_),
    .Y(_0871_)
  );
  NOR _1650_ (
    .A(_0471_),
    .B(_0457_),
    .Y(_0872_)
  );
  NOR _1651_ (
    .A(_1090_),
    .B(_1101_),
    .Y(_0873_)
  );
  NAND _1652_ (
    .A(_0471_),
    .B(_0457_),
    .Y(_0874_)
  );
  NOR _1653_ (
    .A(_0872_),
    .B(_0873_),
    .Y(_0875_)
  );
  NAND _1654_ (
    .A(_0871_),
    .B(_0875_),
    .Y(_0876_)
  );
  NOR _1655_ (
    .A(_0871_),
    .B(_0875_),
    .Y(_0877_)
  );
  NOR _1656_ (
    .A(_0492_),
    .B(_0877_),
    .Y(_0878_)
  );
  NAND _1657_ (
    .A(_0876_),
    .B(_0878_),
    .Y(_0879_)
  );
  NAND _1658_ (
    .A(_0870_),
    .B(_0879_),
    .Y(_0880_)
  );
  NOR _1659_ (
    .A(_0859_),
    .B(_0880_),
    .Y(_0881_)
  );
  NAND _1660_ (
    .A(_0850_),
    .B(_0881_),
    .Y(_1210_)
  );
  NOR _1661_ (
    .A(_0457_),
    .B(_0473_),
    .Y(_0882_)
  );
  NAND _1662_ (
    .A(_0457_),
    .B(_0473_),
    .Y(_0883_)
  );
  NOT _1663_ (
    .A(_0883_),
    .Y(_0884_)
  );
  NOR _1664_ (
    .A(_0882_),
    .B(_0884_),
    .Y(_0885_)
  );
  NOR _1665_ (
    .A(_0842_),
    .B(_0845_),
    .Y(_0886_)
  );
  NOR _1666_ (
    .A(_0843_),
    .B(_0886_),
    .Y(_0887_)
  );
  NOR _1667_ (
    .A(_0885_),
    .B(_0887_),
    .Y(_0888_)
  );
  NAND _1668_ (
    .A(_0885_),
    .B(_0887_),
    .Y(_0889_)
  );
  NOT _1669_ (
    .A(_0889_),
    .Y(_0890_)
  );
  NOR _1670_ (
    .A(_0888_),
    .B(_0890_),
    .Y(_0891_)
  );
  NAND _1671_ (
    .A(_1178_),
    .B(_0891_),
    .Y(_0892_)
  );
  NAND _1672_ (
    .A(_0457_),
    .B(_0474_),
    .Y(_0893_)
  );
  NOT _1673_ (
    .A(_0893_),
    .Y(_0894_)
  );
  NOR _1674_ (
    .A(_0457_),
    .B(_0474_),
    .Y(_0895_)
  );
  NOR _1675_ (
    .A(_0894_),
    .B(_0895_),
    .Y(_0896_)
  );
  NAND _1676_ (
    .A(_0851_),
    .B(_0853_),
    .Y(_0897_)
  );
  NAND _1677_ (
    .A(_0854_),
    .B(_0897_),
    .Y(_0898_)
  );
  NAND _1678_ (
    .A(_0896_),
    .B(_0898_),
    .Y(_0899_)
  );
  NOR _1679_ (
    .A(_0896_),
    .B(_0898_),
    .Y(_0900_)
  );
  NAND _1680_ (
    .A(_0498_),
    .B(_0899_),
    .Y(_0901_)
  );
  NOR _1681_ (
    .A(_0900_),
    .B(_0901_),
    .Y(_0902_)
  );
  NAND _1682_ (
    .A(_0836_),
    .B(_0875_),
    .Y(_0903_)
  );
  NAND _1683_ (
    .A(_0830_),
    .B(_0874_),
    .Y(_0904_)
  );
  NOT _1684_ (
    .A(_0904_),
    .Y(_0905_)
  );
  NAND _1685_ (
    .A(_0903_),
    .B(_0905_),
    .Y(_0906_)
  );
  NAND _1686_ (
    .A(_0457_),
    .B(_0458_),
    .Y(_0907_)
  );
  NOT _1687_ (
    .A(_0907_),
    .Y(_0908_)
  );
  NOR _1688_ (
    .A(_0457_),
    .B(_0458_),
    .Y(_0909_)
  );
  NOR _1689_ (
    .A(_0908_),
    .B(_0909_),
    .Y(_0910_)
  );
  NOR _1690_ (
    .A(_0906_),
    .B(_0910_),
    .Y(_0911_)
  );
  NAND _1691_ (
    .A(_0906_),
    .B(_0910_),
    .Y(_0912_)
  );
  NAND _1692_ (
    .A(_0491_),
    .B(_0912_),
    .Y(_0913_)
  );
  NOR _1693_ (
    .A(_0911_),
    .B(_0913_),
    .Y(_0914_)
  );
  NOR _1694_ (
    .A(_0457_),
    .B(_0862_),
    .Y(_0915_)
  );
  NAND _1695_ (
    .A(_0818_),
    .B(_0873_),
    .Y(_0916_)
  );
  NAND _1696_ (
    .A(_0538_),
    .B(_0916_),
    .Y(_0917_)
  );
  NOR _1697_ (
    .A(_0915_),
    .B(_0917_),
    .Y(_0918_)
  );
  NOR _1698_ (
    .A(_0457_),
    .B(_0535_),
    .Y(_0919_)
  );
  NOR _1699_ (
    .A(_1191_),
    .B(_0882_),
    .Y(_0920_)
  );
  NOR _1700_ (
    .A(_0919_),
    .B(_0920_),
    .Y(_0921_)
  );
  NOR _1701_ (
    .A(_1183_),
    .B(_0883_),
    .Y(_0922_)
  );
  NOR _1702_ (
    .A(_0918_),
    .B(_0922_),
    .Y(_0923_)
  );
  NAND _1703_ (
    .A(_0921_),
    .B(_0923_),
    .Y(_0924_)
  );
  NOR _1704_ (
    .A(_0914_),
    .B(_0924_),
    .Y(_0925_)
  );
  NOT _1705_ (
    .A(_0925_),
    .Y(_0926_)
  );
  NOR _1706_ (
    .A(_0902_),
    .B(_0926_),
    .Y(_0927_)
  );
  NAND _1707_ (
    .A(_0892_),
    .B(_0927_),
    .Y(_1197_)
  );
  NAND _1708_ (
    .A(_0883_),
    .B(_0889_),
    .Y(_0929_)
  );
  NOR _1709_ (
    .A(_0458_),
    .B(_0474_),
    .Y(_0930_)
  );
  NAND _1710_ (
    .A(_0458_),
    .B(_0474_),
    .Y(_0931_)
  );
  NOT _1711_ (
    .A(_0931_),
    .Y(_0932_)
  );
  NOR _1712_ (
    .A(_0930_),
    .B(_0932_),
    .Y(_0933_)
  );
  NAND _1713_ (
    .A(_0929_),
    .B(_0933_),
    .Y(_0934_)
  );
  NOR _1714_ (
    .A(_0929_),
    .B(_0933_),
    .Y(_0935_)
  );
  NOR _1715_ (
    .A(_1179_),
    .B(_0935_),
    .Y(_0936_)
  );
  NAND _1716_ (
    .A(_0934_),
    .B(_0936_),
    .Y(_0937_)
  );
  NAND _1717_ (
    .A(_0893_),
    .B(_0899_),
    .Y(_0938_)
  );
  NOR _1718_ (
    .A(_0458_),
    .B(_0475_),
    .Y(_0940_)
  );
  NAND _1719_ (
    .A(_0458_),
    .B(_0475_),
    .Y(_0941_)
  );
  NOT _1720_ (
    .A(_0941_),
    .Y(_0942_)
  );
  NOR _1721_ (
    .A(_0940_),
    .B(_0942_),
    .Y(_0943_)
  );
  NAND _1722_ (
    .A(_0938_),
    .B(_0943_),
    .Y(_0944_)
  );
  NOR _1723_ (
    .A(_0938_),
    .B(_0943_),
    .Y(_0945_)
  );
  NAND _1724_ (
    .A(_0498_),
    .B(_0944_),
    .Y(_0946_)
  );
  NOR _1725_ (
    .A(_0945_),
    .B(_0946_),
    .Y(_0947_)
  );
  NAND _1726_ (
    .A(_0907_),
    .B(_0912_),
    .Y(_0948_)
  );
  NOR _1727_ (
    .A(_0458_),
    .B(_0459_),
    .Y(_0949_)
  );
  NAND _1728_ (
    .A(_0458_),
    .B(_0459_),
    .Y(_0951_)
  );
  NOT _1729_ (
    .A(_0951_),
    .Y(_0952_)
  );
  NOR _1730_ (
    .A(_0949_),
    .B(_0952_),
    .Y(_0953_)
  );
  NAND _1731_ (
    .A(_0948_),
    .B(_0953_),
    .Y(_0954_)
  );
  NOR _1732_ (
    .A(_0948_),
    .B(_0953_),
    .Y(_0955_)
  );
  NOR _1733_ (
    .A(_0492_),
    .B(_0955_),
    .Y(_0956_)
  );
  NAND _1734_ (
    .A(_0954_),
    .B(_0956_),
    .Y(_0957_)
  );
  NAND _1735_ (
    .A(_1122_),
    .B(_0916_),
    .Y(_0958_)
  );
  NOR _1736_ (
    .A(_0861_),
    .B(_0907_),
    .Y(_0959_)
  );
  NOR _1737_ (
    .A(_0539_),
    .B(_0959_),
    .Y(_0960_)
  );
  NAND _1738_ (
    .A(_0958_),
    .B(_0960_),
    .Y(_0962_)
  );
  NOR _1739_ (
    .A(_0458_),
    .B(_0535_),
    .Y(_0963_)
  );
  NOR _1740_ (
    .A(_1183_),
    .B(_0931_),
    .Y(_0964_)
  );
  NOR _1741_ (
    .A(_1191_),
    .B(_0930_),
    .Y(_0965_)
  );
  NOR _1742_ (
    .A(_0963_),
    .B(_0965_),
    .Y(_0966_)
  );
  NAND _1743_ (
    .A(_0962_),
    .B(_0966_),
    .Y(_0967_)
  );
  NOR _1744_ (
    .A(_0964_),
    .B(_0967_),
    .Y(_0968_)
  );
  NAND _1745_ (
    .A(_0957_),
    .B(_0968_),
    .Y(_0969_)
  );
  NOR _1746_ (
    .A(_0947_),
    .B(_0969_),
    .Y(_0970_)
  );
  NAND _1747_ (
    .A(_0937_),
    .B(_0970_),
    .Y(_1198_)
  );
  NAND _1748_ (
    .A(_0459_),
    .B(_0475_),
    .Y(_0972_)
  );
  NOT _1749_ (
    .A(_0972_),
    .Y(_0973_)
  );
  NOR _1750_ (
    .A(_0459_),
    .B(_0475_),
    .Y(_0974_)
  );
  NOR _1751_ (
    .A(_0973_),
    .B(_0974_),
    .Y(_0975_)
  );
  NOR _1752_ (
    .A(_0929_),
    .B(_0932_),
    .Y(_0976_)
  );
  NOR _1753_ (
    .A(_0930_),
    .B(_0976_),
    .Y(_0977_)
  );
  NAND _1754_ (
    .A(_0975_),
    .B(_0977_),
    .Y(_0978_)
  );
  NOR _1755_ (
    .A(_0975_),
    .B(_0977_),
    .Y(_0979_)
  );
  NOR _1756_ (
    .A(_1179_),
    .B(_0979_),
    .Y(_0980_)
  );
  NAND _1757_ (
    .A(_0978_),
    .B(_0980_),
    .Y(_0981_)
  );
  NAND _1758_ (
    .A(_0459_),
    .B(_0476_),
    .Y(_0983_)
  );
  NOT _1759_ (
    .A(_0983_),
    .Y(_0984_)
  );
  NOR _1760_ (
    .A(_0459_),
    .B(_0476_),
    .Y(_0985_)
  );
  NOR _1761_ (
    .A(_0984_),
    .B(_0985_),
    .Y(_0986_)
  );
  NOR _1762_ (
    .A(_0938_),
    .B(_0942_),
    .Y(_0987_)
  );
  NOR _1763_ (
    .A(_0940_),
    .B(_0987_),
    .Y(_0988_)
  );
  NOR _1764_ (
    .A(_0986_),
    .B(_0988_),
    .Y(_0989_)
  );
  NAND _1765_ (
    .A(_0986_),
    .B(_0988_),
    .Y(_0990_)
  );
  NAND _1766_ (
    .A(_0498_),
    .B(_0990_),
    .Y(_0991_)
  );
  NOR _1767_ (
    .A(_0989_),
    .B(_0991_),
    .Y(_0992_)
  );
  NAND _1768_ (
    .A(_0910_),
    .B(_0953_),
    .Y(_0994_)
  );
  NOT _1769_ (
    .A(_0994_),
    .Y(_0995_)
  );
  NOR _1770_ (
    .A(_0903_),
    .B(_0994_),
    .Y(_0996_)
  );
  NAND _1771_ (
    .A(_0904_),
    .B(_0995_),
    .Y(_0997_)
  );
  NAND _1772_ (
    .A(_0907_),
    .B(_0997_),
    .Y(_0998_)
  );
  NOR _1773_ (
    .A(_0996_),
    .B(_0998_),
    .Y(_0999_)
  );
  NAND _1774_ (
    .A(_0951_),
    .B(_0999_),
    .Y(_1000_)
  );
  NOR _1775_ (
    .A(_0459_),
    .B(_0460_),
    .Y(_1001_)
  );
  NAND _1776_ (
    .A(_0459_),
    .B(_0460_),
    .Y(_1002_)
  );
  NOT _1777_ (
    .A(_1002_),
    .Y(_1003_)
  );
  NOR _1778_ (
    .A(_1001_),
    .B(_1003_),
    .Y(_1005_)
  );
  NAND _1779_ (
    .A(_1000_),
    .B(_1005_),
    .Y(_1006_)
  );
  NOR _1780_ (
    .A(_1000_),
    .B(_1005_),
    .Y(_1007_)
  );
  NOR _1781_ (
    .A(_0492_),
    .B(_1007_),
    .Y(_1008_)
  );
  NAND _1782_ (
    .A(_1006_),
    .B(_1008_),
    .Y(_1009_)
  );
  NOR _1783_ (
    .A(_0459_),
    .B(_0959_),
    .Y(_1010_)
  );
  NOR _1784_ (
    .A(_0916_),
    .B(_0951_),
    .Y(_1011_)
  );
  NOT _1785_ (
    .A(_1011_),
    .Y(_1012_)
  );
  NAND _1786_ (
    .A(_0538_),
    .B(_1012_),
    .Y(_1013_)
  );
  NOR _1787_ (
    .A(_1010_),
    .B(_1013_),
    .Y(_1014_)
  );
  NOR _1788_ (
    .A(_1191_),
    .B(_0974_),
    .Y(_1016_)
  );
  NOR _1789_ (
    .A(_0459_),
    .B(_0535_),
    .Y(_1017_)
  );
  NAND _1790_ (
    .A(_1182_),
    .B(_0973_),
    .Y(_1018_)
  );
  NOR _1791_ (
    .A(_1016_),
    .B(_1017_),
    .Y(_1019_)
  );
  NAND _1792_ (
    .A(_1018_),
    .B(_1019_),
    .Y(_1020_)
  );
  NOR _1793_ (
    .A(_1014_),
    .B(_1020_),
    .Y(_1021_)
  );
  NAND _1794_ (
    .A(_1009_),
    .B(_1021_),
    .Y(_1022_)
  );
  NOR _1795_ (
    .A(_0992_),
    .B(_1022_),
    .Y(_1023_)
  );
  NAND _1796_ (
    .A(_0981_),
    .B(_1023_),
    .Y(_1199_)
  );
  NAND _1797_ (
    .A(_0972_),
    .B(_0978_),
    .Y(_1024_)
  );
  NAND _1798_ (
    .A(_0460_),
    .B(_0476_),
    .Y(_1026_)
  );
  NOR _1799_ (
    .A(_0460_),
    .B(_0476_),
    .Y(_1027_)
  );
  NAND _1800_ (
    .A(_1133_),
    .B(_1144_),
    .Y(_1028_)
  );
  NAND _1801_ (
    .A(_1026_),
    .B(_1028_),
    .Y(_1029_)
  );
  NAND _1802_ (
    .A(_1024_),
    .B(_1029_),
    .Y(_1030_)
  );
  NOT _1803_ (
    .A(_1030_),
    .Y(_1031_)
  );
  NOR _1804_ (
    .A(_1024_),
    .B(_1029_),
    .Y(_1032_)
  );
  NOR _1805_ (
    .A(_1031_),
    .B(_1032_),
    .Y(_1033_)
  );
  NOR _1806_ (
    .A(_1179_),
    .B(_1033_),
    .Y(_1034_)
  );
  NAND _1807_ (
    .A(_0983_),
    .B(_0990_),
    .Y(_1035_)
  );
  NOR _1808_ (
    .A(_0460_),
    .B(_0477_),
    .Y(_1037_)
  );
  NAND _1809_ (
    .A(_0460_),
    .B(_0477_),
    .Y(_1038_)
  );
  NOT _1810_ (
    .A(_1038_),
    .Y(_1039_)
  );
  NOR _1811_ (
    .A(_1037_),
    .B(_1039_),
    .Y(_1040_)
  );
  NAND _1812_ (
    .A(_1035_),
    .B(_1040_),
    .Y(_1041_)
  );
  NOR _1813_ (
    .A(_1035_),
    .B(_1040_),
    .Y(_1042_)
  );
  NAND _1814_ (
    .A(_0498_),
    .B(_1041_),
    .Y(_1043_)
  );
  NOR _1815_ (
    .A(_1042_),
    .B(_1043_),
    .Y(_1044_)
  );
  NAND _1816_ (
    .A(_1002_),
    .B(_1006_),
    .Y(_1045_)
  );
  NOR _1817_ (
    .A(_0460_),
    .B(_0461_),
    .Y(_1046_)
  );
  NAND _1818_ (
    .A(_0460_),
    .B(_0461_),
    .Y(_1048_)
  );
  NOT _1819_ (
    .A(_1048_),
    .Y(_1049_)
  );
  NOR _1820_ (
    .A(_1046_),
    .B(_1049_),
    .Y(_1050_)
  );
  NOT _1821_ (
    .A(_1050_),
    .Y(_1051_)
  );
  NAND _1822_ (
    .A(_1045_),
    .B(_1050_),
    .Y(_1052_)
  );
  NOR _1823_ (
    .A(_1045_),
    .B(_1050_),
    .Y(_1053_)
  );
  NOR _1824_ (
    .A(_0492_),
    .B(_1053_),
    .Y(_1054_)
  );
  NAND _1825_ (
    .A(_1052_),
    .B(_1054_),
    .Y(_1055_)
  );
  NOR _1826_ (
    .A(_0460_),
    .B(_1011_),
    .Y(_1056_)
  );
  NOR _1827_ (
    .A(_1133_),
    .B(_1012_),
    .Y(_1057_)
  );
  NAND _1828_ (
    .A(_0460_),
    .B(_1011_),
    .Y(_1059_)
  );
  NOR _1829_ (
    .A(_1056_),
    .B(_1057_),
    .Y(_1060_)
  );
  NAND _1830_ (
    .A(_0538_),
    .B(_1060_),
    .Y(_1061_)
  );
  NOR _1831_ (
    .A(_1183_),
    .B(_1026_),
    .Y(_1062_)
  );
  NOR _1832_ (
    .A(_1191_),
    .B(_1027_),
    .Y(_1063_)
  );
  NOR _1833_ (
    .A(_0460_),
    .B(_0535_),
    .Y(_1064_)
  );
  NOR _1834_ (
    .A(_1063_),
    .B(_1064_),
    .Y(_1065_)
  );
  NAND _1835_ (
    .A(_1061_),
    .B(_1065_),
    .Y(_1066_)
  );
  NOR _1836_ (
    .A(_1062_),
    .B(_1066_),
    .Y(_1067_)
  );
  NAND _1837_ (
    .A(_1055_),
    .B(_1067_),
    .Y(_1068_)
  );
  NOR _1838_ (
    .A(_1044_),
    .B(_1068_),
    .Y(_1070_)
  );
  NOT _1839_ (
    .A(_1070_),
    .Y(_1071_)
  );
  NOR _1840_ (
    .A(_1034_),
    .B(_1071_),
    .Y(_1072_)
  );
  NOT _1841_ (
    .A(_1072_),
    .Y(_1200_)
  );
  NAND _1842_ (
    .A(_0461_),
    .B(_0477_),
    .Y(_1073_)
  );
  NOT _1843_ (
    .A(_1073_),
    .Y(_1074_)
  );
  NOR _1844_ (
    .A(_0461_),
    .B(_0477_),
    .Y(_1075_)
  );
  NOR _1845_ (
    .A(_1074_),
    .B(_1075_),
    .Y(_1076_)
  );
  NAND _1846_ (
    .A(_1024_),
    .B(_1028_),
    .Y(_1077_)
  );
  NAND _1847_ (
    .A(_1026_),
    .B(_1077_),
    .Y(_1078_)
  );
  NAND _1848_ (
    .A(_1076_),
    .B(_1078_),
    .Y(_1080_)
  );
  NOR _1849_ (
    .A(_1076_),
    .B(_1078_),
    .Y(_1081_)
  );
  NOR _1850_ (
    .A(_1179_),
    .B(_1081_),
    .Y(_1082_)
  );
  NAND _1851_ (
    .A(_1080_),
    .B(_1082_),
    .Y(_1083_)
  );
  NOR _1852_ (
    .A(_0461_),
    .B(_0478_),
    .Y(_1084_)
  );
  NAND _1853_ (
    .A(_0461_),
    .B(_0478_),
    .Y(_1085_)
  );
  NOT _1854_ (
    .A(_1085_),
    .Y(_1086_)
  );
  NOR _1855_ (
    .A(_1084_),
    .B(_1086_),
    .Y(_1087_)
  );
  NOR _1856_ (
    .A(_1035_),
    .B(_1039_),
    .Y(_1088_)
  );
  NOR _1857_ (
    .A(_1037_),
    .B(_1088_),
    .Y(_1089_)
  );
  NAND _1858_ (
    .A(_1087_),
    .B(_1089_),
    .Y(_1091_)
  );
  NOR _1859_ (
    .A(_1087_),
    .B(_1089_),
    .Y(_1092_)
  );
  NAND _1860_ (
    .A(_0498_),
    .B(_1091_),
    .Y(_1093_)
  );
  NOR _1861_ (
    .A(_1092_),
    .B(_1093_),
    .Y(_1094_)
  );
  NOR _1862_ (
    .A(_1006_),
    .B(_1051_),
    .Y(_1095_)
  );
  NAND _1863_ (
    .A(_1002_),
    .B(_1048_),
    .Y(_1096_)
  );
  NOR _1864_ (
    .A(_1095_),
    .B(_1096_),
    .Y(_1097_)
  );
  NOT _1865_ (
    .A(_1097_),
    .Y(_1098_)
  );
  NOR _1866_ (
    .A(_0461_),
    .B(_1165_),
    .Y(_1099_)
  );
  NOR _1867_ (
    .A(_1154_),
    .B(_0462_),
    .Y(_1100_)
  );
  NOR _1868_ (
    .A(_1099_),
    .B(_1100_),
    .Y(_1102_)
  );
  NAND _1869_ (
    .A(_1097_),
    .B(_1102_),
    .Y(_1103_)
  );
  NOR _1870_ (
    .A(_1097_),
    .B(_1102_),
    .Y(_1104_)
  );
  NOR _1871_ (
    .A(_0492_),
    .B(_1104_),
    .Y(_1105_)
  );
  NAND _1872_ (
    .A(_1103_),
    .B(_1105_),
    .Y(_1106_)
  );
  NAND _1873_ (
    .A(_1154_),
    .B(_1059_),
    .Y(_1107_)
  );
  NAND _1874_ (
    .A(_0461_),
    .B(_1057_),
    .Y(_1108_)
  );
  NAND _1875_ (
    .A(_0950_),
    .B(_1108_),
    .Y(_1109_)
  );
  NOR _1876_ (
    .A(_1186_),
    .B(_1109_),
    .Y(_1110_)
  );
  NAND _1877_ (
    .A(_1107_),
    .B(_1110_),
    .Y(_1111_)
  );
  NOR _1878_ (
    .A(_1191_),
    .B(_1075_),
    .Y(_1113_)
  );
  NOR _1879_ (
    .A(_1183_),
    .B(_1073_),
    .Y(_1114_)
  );
  NOR _1880_ (
    .A(_0461_),
    .B(_0535_),
    .Y(_1115_)
  );
  NOR _1881_ (
    .A(_1113_),
    .B(_1114_),
    .Y(_1116_)
  );
  NAND _1882_ (
    .A(_1111_),
    .B(_1116_),
    .Y(_1117_)
  );
  NOR _1883_ (
    .A(_1115_),
    .B(_1117_),
    .Y(_1118_)
  );
  NAND _1884_ (
    .A(_1106_),
    .B(_1118_),
    .Y(_1119_)
  );
  NOR _1885_ (
    .A(_1094_),
    .B(_1119_),
    .Y(_1120_)
  );
  NAND _1886_ (
    .A(_1083_),
    .B(_1120_),
    .Y(_1201_)
  );
  NAND _1887_ (
    .A(_1073_),
    .B(_1080_),
    .Y(_1121_)
  );
  NOR _1888_ (
    .A(_0462_),
    .B(_0478_),
    .Y(_1123_)
  );
  NAND _1889_ (
    .A(_0462_),
    .B(_0478_),
    .Y(_1124_)
  );
  NOT _1890_ (
    .A(_1124_),
    .Y(_1125_)
  );
  NOR _1891_ (
    .A(_1123_),
    .B(_1125_),
    .Y(_1126_)
  );
  NOR _1892_ (
    .A(_1121_),
    .B(_1126_),
    .Y(_1127_)
  );
  NAND _1893_ (
    .A(_1121_),
    .B(_1126_),
    .Y(_1128_)
  );
  NOR _1894_ (
    .A(_1179_),
    .B(_1127_),
    .Y(_1129_)
  );
  NAND _1895_ (
    .A(_1128_),
    .B(_1129_),
    .Y(_1130_)
  );
  NAND _1896_ (
    .A(_1085_),
    .B(_1091_),
    .Y(_1131_)
  );
  NAND _1897_ (
    .A(_0462_),
    .B(_1131_),
    .Y(_1132_)
  );
  NOR _1898_ (
    .A(_0462_),
    .B(_1131_),
    .Y(_1134_)
  );
  NAND _1899_ (
    .A(_0498_),
    .B(_1132_),
    .Y(_1135_)
  );
  NOR _1900_ (
    .A(_1134_),
    .B(_1135_),
    .Y(_1136_)
  );
  NOR _1901_ (
    .A(_1099_),
    .B(_1104_),
    .Y(_1137_)
  );
  NAND _1902_ (
    .A(_1098_),
    .B(_1099_),
    .Y(_1138_)
  );
  NAND _1903_ (
    .A(_0491_),
    .B(_1138_),
    .Y(_1139_)
  );
  NOR _1904_ (
    .A(_1137_),
    .B(_1139_),
    .Y(_1140_)
  );
  NAND _1905_ (
    .A(_0462_),
    .B(_1110_),
    .Y(_1141_)
  );
  NOR _1906_ (
    .A(_0462_),
    .B(_1186_),
    .Y(_1142_)
  );
  NAND _1907_ (
    .A(_1109_),
    .B(_1142_),
    .Y(_1143_)
  );
  NOR _1908_ (
    .A(_1191_),
    .B(_1123_),
    .Y(_1145_)
  );
  NOR _1909_ (
    .A(_1183_),
    .B(_1124_),
    .Y(_1146_)
  );
  NOR _1910_ (
    .A(_1145_),
    .B(_1146_),
    .Y(_1147_)
  );
  NAND _1911_ (
    .A(_1141_),
    .B(_1147_),
    .Y(_1148_)
  );
  NOR _1912_ (
    .A(_1140_),
    .B(_1148_),
    .Y(_1149_)
  );
  NAND _1913_ (
    .A(_1143_),
    .B(_1149_),
    .Y(_1150_)
  );
  NOR _1914_ (
    .A(_1136_),
    .B(_1150_),
    .Y(_1151_)
  );
  NAND _1915_ (
    .A(_1130_),
    .B(_1151_),
    .Y(_0488_)
  );
  NOR _1916_ (
    .A(_1198_),
    .B(_1201_),
    .Y(_1152_)
  );
  NOR _1917_ (
    .A(_1206_),
    .B(_1207_),
    .Y(_1153_)
  );
  NAND _1918_ (
    .A(_0507_),
    .B(_1153_),
    .Y(_1155_)
  );
  NOR _1919_ (
    .A(_1199_),
    .B(_1155_),
    .Y(_1156_)
  );
  NOT _1920_ (
    .A(_1156_),
    .Y(_1157_)
  );
  NOR _1921_ (
    .A(_1204_),
    .B(_1208_),
    .Y(_1158_)
  );
  NOT _1922_ (
    .A(_1158_),
    .Y(_1159_)
  );
  NOR _1923_ (
    .A(_1205_),
    .B(_1159_),
    .Y(_1160_)
  );
  NOR _1924_ (
    .A(_1209_),
    .B(_1210_),
    .Y(_1161_)
  );
  NAND _1925_ (
    .A(_1160_),
    .B(_1161_),
    .Y(_1162_)
  );
  NOR _1926_ (
    .A(_1157_),
    .B(_1162_),
    .Y(_1163_)
  );
  NAND _1927_ (
    .A(_1072_),
    .B(_1163_),
    .Y(_1164_)
  );
  NOR _1928_ (
    .A(_1203_),
    .B(_1197_),
    .Y(_1166_)
  );
  NAND _1929_ (
    .A(_0546_),
    .B(_1166_),
    .Y(_1167_)
  );
  NOR _1930_ (
    .A(_1164_),
    .B(_1167_),
    .Y(_1168_)
  );
  NAND _1931_ (
    .A(_1152_),
    .B(_1168_),
    .Y(_1169_)
  );
  NOR _1932_ (
    .A(_0488_),
    .B(_1169_),
    .Y(_1211_)
  );
  assign outF[15] = neg;
  assign _1193_ = opc[0];
  assign _1194_ = opc[1];
  assign _1195_ = opc[2];
  assign _0472_ = inN[0];
  assign _0456_ = inM[0];
  assign _0463_ = inM[1];
  assign _0479_ = inN[1];
  assign _0455_ = inC;
  assign outF[0] = _1196_;
  assign _0464_ = inM[2];
  assign _0480_ = inN[2];
  assign outF[1] = _1202_;
  assign _0465_ = inM[3];
  assign _0481_ = inN[3];
  assign outF[2] = _1203_;
  assign _0466_ = inM[4];
  assign _0482_ = inN[4];
  assign outF[3] = _1204_;
  assign _0467_ = inM[5];
  assign _0483_ = inN[5];
  assign outF[4] = _1205_;
  assign _0468_ = inM[6];
  assign _0484_ = inN[6];
  assign outF[5] = _1206_;
  assign _0469_ = inM[7];
  assign _0485_ = inN[7];
  assign outF[6] = _1207_;
  assign _0470_ = inM[8];
  assign _0486_ = inN[8];
  assign outF[7] = _1208_;
  assign _0471_ = inM[9];
  assign _0487_ = inN[9];
  assign outF[8] = _1209_;
  assign _0457_ = inM[10];
  assign _0473_ = inN[10];
  assign outF[9] = _1210_;
  assign _0458_ = inM[11];
  assign _0474_ = inN[11];
  assign outF[10] = _1197_;
  assign _0459_ = inM[12];
  assign _0475_ = inN[12];
  assign outF[11] = _1198_;
  assign _0460_ = inM[13];
  assign _0476_ = inN[13];
  assign outF[12] = _1199_;
  assign _0461_ = inM[14];
  assign _0477_ = inN[14];
  assign outF[13] = _1200_;
  assign _0462_ = inM[15];
  assign _0478_ = inN[15];
  assign outF[14] = _1201_;
  assign neg = _0488_;
  assign zer = _1211_;
endmodule
