`timescale 1ns/1ns
module Q2 (input signed [15:0] inM, inN, input inC, input [2:0] opc, output signed [15:0] outF, output zer, neg);
	wire [15:0] wAdd, wAnd, wOr, wInv, wShif1, wShif2, wMux;
	wire w1, w2, w3, w4, w5, w6, co;
	assign neg = outF[15];
	Shifter2bit1 S1(inN, wShif1);
	Shifter2bit1 S2(inM, wShif2);
	or O1(w1, opc[1], opc[0]);
	not N1(w2, opc[2]);
	not N2(zer, w5);
	and A2(w3, opc[2], w1);
	and A3(w4, opc[0], w2);
	nor N3(w6, opc[0], opc[1], opc[2]);
	Mux4 M1(wAdd, wAnd, wOr, wInv, {w3,w4}, outF);
	Mux4 M2(inN, wShif1, 16'b1, wShif2, {opc[1], opc[0]}, wMux);
	Orbits G4(outF, w5);
	Adder A1(inM, wMux, w6, co, wAdd);
	Inventer G1(inM, wInv);
	And16bit G3(inM, inN, wAnd);
	Or16bit G2(inM, inN, wOr);
endmodule

module Shifter2bit1 (input signed [15:0] A, output signed [15:0] W);
	assign W = A >>> 1;
endmodule

module Adder (input signed [15:0] A,B, input ci, output signed [15:0] W, output co);
	assign {co,W}= A + B + ci;
endmodule

module And16bit (input [15:0] A,B, output [15:0] W);
	assign W = A & B;
endmodule

module Mux4 (input [15:0] A1, A2, A3, A4,input [1:0] select,output [15:0] W);
	assign W =	(select==2'd0) ? A1:
			(select==2'd1) ? A2:
			(select==2'd2) ? A3:
			(select==2'd3) ? A4:
			16'bx;
endmodule

module Mux2 (input A1, A2,select,output W);
	assign W =	(select==1'b0) ? A1: 
			(select==1'b1) ? A2:
			1'bx;
endmodule

module Or16bit (input [15:0] A,B, output [15:0] W);
	assign W = A | B;
endmodule

module Orbits (input [15:0] A, output W);
	assign W = | A;
endmodule

module Inventer (input [15:0] A, output [15:0] W);
	assign W = ~ A;
endmodule

module NOT(A, Y);
input A;
output Y;
assign Y = ~A;
endmodule

module NAND(A, B, Y);
input A, B;
output Y;
assign Y = ~(A & B);
endmodule

module NOR(A, B, Y);
input A, B;
output Y;
assign Y = ~(A | B);
endmodule

module DFF(C, D, Q);
input C, D;
output reg Q;
always @(posedge C)
	Q <= D;
endmodule

module Adder(A, B, ci, W, co);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire _272_;
  wire _273_;
  wire _274_;
  wire _275_;
  wire _276_;
  wire _277_;
  wire _278_;
  wire _279_;
  wire _280_;
  wire _281_;
  wire _282_;
  wire _283_;
  wire _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire _304_;
  wire _305_;
  wire _306_;
  wire _307_;
  wire _308_;
  wire _309_;
  wire _310_;
  wire _311_;
  wire _312_;
  wire _313_;
  wire _314_;
  wire _315_;
  wire _316_;
  wire _317_;
  wire _318_;
  wire _319_;
  wire _320_;
  wire _321_;
  wire _322_;
  wire _323_;
  wire _324_;
  wire _325_;
  wire _326_;
  wire _327_;
  wire _328_;
  wire _329_;
  wire _330_;
  wire _331_;
  wire _332_;
  wire _333_;
  wire _334_;
  input [15:0] A;
  input [15:0] B;
  output [15:0] W;
  input ci;
  output co;
  NOT _335_ (
    .A(_098_),
    .Y(_287_)
  );
  NOT _336_ (
    .A(_082_),
    .Y(_288_)
  );
  NOT _337_ (
    .A(_130_),
    .Y(_289_)
  );
  NOT _338_ (
    .A(_105_),
    .Y(_290_)
  );
  NOT _339_ (
    .A(_089_),
    .Y(_291_)
  );
  NOT _340_ (
    .A(_106_),
    .Y(_292_)
  );
  NOT _341_ (
    .A(_090_),
    .Y(_293_)
  );
  NOT _342_ (
    .A(_107_),
    .Y(_294_)
  );
  NOT _343_ (
    .A(_091_),
    .Y(_295_)
  );
  NOT _344_ (
    .A(_108_),
    .Y(_296_)
  );
  NOT _345_ (
    .A(_092_),
    .Y(_297_)
  );
  NOT _346_ (
    .A(_109_),
    .Y(_298_)
  );
  NOT _347_ (
    .A(_093_),
    .Y(_299_)
  );
  NOT _348_ (
    .A(_110_),
    .Y(_300_)
  );
  NOT _349_ (
    .A(_094_),
    .Y(_301_)
  );
  NOT _350_ (
    .A(_111_),
    .Y(_302_)
  );
  NOT _351_ (
    .A(_095_),
    .Y(_303_)
  );
  NOT _352_ (
    .A(_112_),
    .Y(_304_)
  );
  NOT _353_ (
    .A(_096_),
    .Y(_305_)
  );
  NOT _354_ (
    .A(_113_),
    .Y(_306_)
  );
  NOT _355_ (
    .A(_097_),
    .Y(_307_)
  );
  NOT _356_ (
    .A(_099_),
    .Y(_308_)
  );
  NOT _357_ (
    .A(_083_),
    .Y(_309_)
  );
  NOT _358_ (
    .A(_100_),
    .Y(_310_)
  );
  NOT _359_ (
    .A(_084_),
    .Y(_311_)
  );
  NOT _360_ (
    .A(_101_),
    .Y(_312_)
  );
  NOT _361_ (
    .A(_085_),
    .Y(_313_)
  );
  NOT _362_ (
    .A(_102_),
    .Y(_314_)
  );
  NOT _363_ (
    .A(_086_),
    .Y(_315_)
  );
  NOT _364_ (
    .A(_103_),
    .Y(_316_)
  );
  NOT _365_ (
    .A(_087_),
    .Y(_317_)
  );
  NOT _366_ (
    .A(_104_),
    .Y(_318_)
  );
  NOT _367_ (
    .A(_088_),
    .Y(_319_)
  );
  NOR _368_ (
    .A(_287_),
    .B(_288_),
    .Y(_320_)
  );
  NAND _369_ (
    .A(_098_),
    .B(_082_),
    .Y(_321_)
  );
  NOR _370_ (
    .A(_098_),
    .B(_082_),
    .Y(_322_)
  );
  NOT _371_ (
    .A(_322_),
    .Y(_323_)
  );
  NOR _372_ (
    .A(_320_),
    .B(_322_),
    .Y(_324_)
  );
  NAND _373_ (
    .A(_321_),
    .B(_323_),
    .Y(_325_)
  );
  NOR _374_ (
    .A(_289_),
    .B(_325_),
    .Y(_326_)
  );
  NAND _375_ (
    .A(_130_),
    .B(_324_),
    .Y(_327_)
  );
  NOR _376_ (
    .A(_130_),
    .B(_324_),
    .Y(_328_)
  );
  NOR _377_ (
    .A(_326_),
    .B(_328_),
    .Y(_114_)
  );
  NOR _378_ (
    .A(_320_),
    .B(_326_),
    .Y(_329_)
  );
  NAND _379_ (
    .A(_321_),
    .B(_327_),
    .Y(_330_)
  );
  NOR _380_ (
    .A(_105_),
    .B(_089_),
    .Y(_331_)
  );
  NOR _381_ (
    .A(_290_),
    .B(_291_),
    .Y(_332_)
  );
  NAND _382_ (
    .A(_105_),
    .B(_089_),
    .Y(_333_)
  );
  NOR _383_ (
    .A(_331_),
    .B(_332_),
    .Y(_334_)
  );
  NOT _384_ (
    .A(_334_),
    .Y(_132_)
  );
  NOR _385_ (
    .A(_329_),
    .B(_132_),
    .Y(_133_)
  );
  NAND _386_ (
    .A(_330_),
    .B(_334_),
    .Y(_134_)
  );
  NOR _387_ (
    .A(_330_),
    .B(_334_),
    .Y(_135_)
  );
  NOR _388_ (
    .A(_133_),
    .B(_135_),
    .Y(_121_)
  );
  NOR _389_ (
    .A(_332_),
    .B(_133_),
    .Y(_136_)
  );
  NAND _390_ (
    .A(_333_),
    .B(_134_),
    .Y(_137_)
  );
  NOR _391_ (
    .A(_106_),
    .B(_090_),
    .Y(_138_)
  );
  NOR _392_ (
    .A(_292_),
    .B(_293_),
    .Y(_139_)
  );
  NAND _393_ (
    .A(_106_),
    .B(_090_),
    .Y(_140_)
  );
  NOR _394_ (
    .A(_138_),
    .B(_139_),
    .Y(_141_)
  );
  NOT _395_ (
    .A(_141_),
    .Y(_142_)
  );
  NOR _396_ (
    .A(_136_),
    .B(_142_),
    .Y(_143_)
  );
  NAND _397_ (
    .A(_137_),
    .B(_141_),
    .Y(_144_)
  );
  NOR _398_ (
    .A(_137_),
    .B(_141_),
    .Y(_145_)
  );
  NOR _399_ (
    .A(_143_),
    .B(_145_),
    .Y(_122_)
  );
  NOR _400_ (
    .A(_139_),
    .B(_143_),
    .Y(_146_)
  );
  NAND _401_ (
    .A(_140_),
    .B(_144_),
    .Y(_147_)
  );
  NOR _402_ (
    .A(_107_),
    .B(_091_),
    .Y(_148_)
  );
  NAND _403_ (
    .A(_294_),
    .B(_295_),
    .Y(_149_)
  );
  NOR _404_ (
    .A(_294_),
    .B(_295_),
    .Y(_150_)
  );
  NAND _405_ (
    .A(_107_),
    .B(_091_),
    .Y(_151_)
  );
  NOR _406_ (
    .A(_148_),
    .B(_150_),
    .Y(_152_)
  );
  NAND _407_ (
    .A(_149_),
    .B(_151_),
    .Y(_153_)
  );
  NAND _408_ (
    .A(_146_),
    .B(_152_),
    .Y(_154_)
  );
  NAND _409_ (
    .A(_147_),
    .B(_153_),
    .Y(_155_)
  );
  NAND _410_ (
    .A(_154_),
    .B(_155_),
    .Y(_123_)
  );
  NOR _411_ (
    .A(_296_),
    .B(_297_),
    .Y(_156_)
  );
  NAND _412_ (
    .A(_108_),
    .B(_092_),
    .Y(_157_)
  );
  NOR _413_ (
    .A(_108_),
    .B(_092_),
    .Y(_158_)
  );
  NOR _414_ (
    .A(_156_),
    .B(_158_),
    .Y(_159_)
  );
  NOT _415_ (
    .A(_159_),
    .Y(_160_)
  );
  NOR _416_ (
    .A(_146_),
    .B(_148_),
    .Y(_161_)
  );
  NAND _417_ (
    .A(_147_),
    .B(_149_),
    .Y(_162_)
  );
  NOR _418_ (
    .A(_150_),
    .B(_161_),
    .Y(_163_)
  );
  NAND _419_ (
    .A(_151_),
    .B(_162_),
    .Y(_164_)
  );
  NOR _420_ (
    .A(_160_),
    .B(_163_),
    .Y(_165_)
  );
  NAND _421_ (
    .A(_159_),
    .B(_164_),
    .Y(_166_)
  );
  NOR _422_ (
    .A(_159_),
    .B(_164_),
    .Y(_167_)
  );
  NOR _423_ (
    .A(_165_),
    .B(_167_),
    .Y(_124_)
  );
  NOR _424_ (
    .A(_156_),
    .B(_165_),
    .Y(_168_)
  );
  NAND _425_ (
    .A(_157_),
    .B(_166_),
    .Y(_169_)
  );
  NOR _426_ (
    .A(_109_),
    .B(_093_),
    .Y(_170_)
  );
  NOR _427_ (
    .A(_298_),
    .B(_299_),
    .Y(_171_)
  );
  NAND _428_ (
    .A(_109_),
    .B(_093_),
    .Y(_172_)
  );
  NOR _429_ (
    .A(_170_),
    .B(_171_),
    .Y(_173_)
  );
  NOT _430_ (
    .A(_173_),
    .Y(_174_)
  );
  NOR _431_ (
    .A(_168_),
    .B(_174_),
    .Y(_175_)
  );
  NAND _432_ (
    .A(_169_),
    .B(_173_),
    .Y(_176_)
  );
  NOR _433_ (
    .A(_169_),
    .B(_173_),
    .Y(_177_)
  );
  NOR _434_ (
    .A(_175_),
    .B(_177_),
    .Y(_125_)
  );
  NOR _435_ (
    .A(_171_),
    .B(_175_),
    .Y(_178_)
  );
  NAND _436_ (
    .A(_172_),
    .B(_176_),
    .Y(_179_)
  );
  NOR _437_ (
    .A(_110_),
    .B(_094_),
    .Y(_180_)
  );
  NOR _438_ (
    .A(_300_),
    .B(_301_),
    .Y(_181_)
  );
  NAND _439_ (
    .A(_110_),
    .B(_094_),
    .Y(_182_)
  );
  NOR _440_ (
    .A(_180_),
    .B(_181_),
    .Y(_183_)
  );
  NOT _441_ (
    .A(_183_),
    .Y(_184_)
  );
  NOR _442_ (
    .A(_178_),
    .B(_184_),
    .Y(_185_)
  );
  NAND _443_ (
    .A(_179_),
    .B(_183_),
    .Y(_186_)
  );
  NOR _444_ (
    .A(_179_),
    .B(_183_),
    .Y(_187_)
  );
  NOR _445_ (
    .A(_185_),
    .B(_187_),
    .Y(_126_)
  );
  NOR _446_ (
    .A(_181_),
    .B(_185_),
    .Y(_188_)
  );
  NAND _447_ (
    .A(_182_),
    .B(_186_),
    .Y(_189_)
  );
  NOR _448_ (
    .A(_111_),
    .B(_095_),
    .Y(_190_)
  );
  NAND _449_ (
    .A(_302_),
    .B(_303_),
    .Y(_191_)
  );
  NOR _450_ (
    .A(_302_),
    .B(_303_),
    .Y(_192_)
  );
  NAND _451_ (
    .A(_111_),
    .B(_095_),
    .Y(_193_)
  );
  NOR _452_ (
    .A(_190_),
    .B(_192_),
    .Y(_194_)
  );
  NAND _453_ (
    .A(_191_),
    .B(_193_),
    .Y(_195_)
  );
  NOR _454_ (
    .A(_189_),
    .B(_194_),
    .Y(_196_)
  );
  NOR _455_ (
    .A(_188_),
    .B(_195_),
    .Y(_197_)
  );
  NOR _456_ (
    .A(_196_),
    .B(_197_),
    .Y(_127_)
  );
  NOR _457_ (
    .A(_112_),
    .B(_096_),
    .Y(_198_)
  );
  NOR _458_ (
    .A(_304_),
    .B(_305_),
    .Y(_199_)
  );
  NAND _459_ (
    .A(_112_),
    .B(_096_),
    .Y(_200_)
  );
  NOR _460_ (
    .A(_198_),
    .B(_199_),
    .Y(_201_)
  );
  NOT _461_ (
    .A(_201_),
    .Y(_202_)
  );
  NOR _462_ (
    .A(_188_),
    .B(_190_),
    .Y(_203_)
  );
  NAND _463_ (
    .A(_189_),
    .B(_191_),
    .Y(_204_)
  );
  NOR _464_ (
    .A(_192_),
    .B(_203_),
    .Y(_205_)
  );
  NAND _465_ (
    .A(_193_),
    .B(_204_),
    .Y(_206_)
  );
  NOR _466_ (
    .A(_202_),
    .B(_205_),
    .Y(_207_)
  );
  NAND _467_ (
    .A(_201_),
    .B(_206_),
    .Y(_208_)
  );
  NOR _468_ (
    .A(_201_),
    .B(_206_),
    .Y(_209_)
  );
  NOR _469_ (
    .A(_207_),
    .B(_209_),
    .Y(_128_)
  );
  NOR _470_ (
    .A(_199_),
    .B(_207_),
    .Y(_210_)
  );
  NAND _471_ (
    .A(_200_),
    .B(_208_),
    .Y(_211_)
  );
  NOR _472_ (
    .A(_113_),
    .B(_097_),
    .Y(_212_)
  );
  NAND _473_ (
    .A(_306_),
    .B(_307_),
    .Y(_213_)
  );
  NOR _474_ (
    .A(_306_),
    .B(_307_),
    .Y(_214_)
  );
  NAND _475_ (
    .A(_113_),
    .B(_097_),
    .Y(_215_)
  );
  NOR _476_ (
    .A(_212_),
    .B(_214_),
    .Y(_216_)
  );
  NAND _477_ (
    .A(_213_),
    .B(_215_),
    .Y(_217_)
  );
  NAND _478_ (
    .A(_211_),
    .B(_217_),
    .Y(_218_)
  );
  NAND _479_ (
    .A(_210_),
    .B(_216_),
    .Y(_219_)
  );
  NAND _480_ (
    .A(_218_),
    .B(_219_),
    .Y(_129_)
  );
  NOR _481_ (
    .A(_308_),
    .B(_309_),
    .Y(_220_)
  );
  NAND _482_ (
    .A(_099_),
    .B(_083_),
    .Y(_221_)
  );
  NOR _483_ (
    .A(_099_),
    .B(_083_),
    .Y(_222_)
  );
  NOR _484_ (
    .A(_220_),
    .B(_222_),
    .Y(_223_)
  );
  NOT _485_ (
    .A(_223_),
    .Y(_224_)
  );
  NOR _486_ (
    .A(_211_),
    .B(_214_),
    .Y(_225_)
  );
  NAND _487_ (
    .A(_210_),
    .B(_215_),
    .Y(_226_)
  );
  NOR _488_ (
    .A(_212_),
    .B(_225_),
    .Y(_227_)
  );
  NAND _489_ (
    .A(_213_),
    .B(_226_),
    .Y(_228_)
  );
  NOR _490_ (
    .A(_224_),
    .B(_228_),
    .Y(_229_)
  );
  NAND _491_ (
    .A(_223_),
    .B(_227_),
    .Y(_230_)
  );
  NOR _492_ (
    .A(_223_),
    .B(_227_),
    .Y(_231_)
  );
  NOR _493_ (
    .A(_229_),
    .B(_231_),
    .Y(_115_)
  );
  NOR _494_ (
    .A(_220_),
    .B(_229_),
    .Y(_232_)
  );
  NAND _495_ (
    .A(_221_),
    .B(_230_),
    .Y(_233_)
  );
  NOR _496_ (
    .A(_100_),
    .B(_084_),
    .Y(_234_)
  );
  NAND _497_ (
    .A(_310_),
    .B(_311_),
    .Y(_235_)
  );
  NOR _498_ (
    .A(_310_),
    .B(_311_),
    .Y(_236_)
  );
  NAND _499_ (
    .A(_100_),
    .B(_084_),
    .Y(_237_)
  );
  NOR _500_ (
    .A(_234_),
    .B(_236_),
    .Y(_238_)
  );
  NAND _501_ (
    .A(_235_),
    .B(_237_),
    .Y(_239_)
  );
  NAND _502_ (
    .A(_233_),
    .B(_239_),
    .Y(_240_)
  );
  NAND _503_ (
    .A(_232_),
    .B(_238_),
    .Y(_241_)
  );
  NAND _504_ (
    .A(_240_),
    .B(_241_),
    .Y(_116_)
  );
  NOR _505_ (
    .A(_101_),
    .B(_085_),
    .Y(_242_)
  );
  NOR _506_ (
    .A(_312_),
    .B(_313_),
    .Y(_243_)
  );
  NAND _507_ (
    .A(_101_),
    .B(_085_),
    .Y(_244_)
  );
  NOR _508_ (
    .A(_242_),
    .B(_243_),
    .Y(_245_)
  );
  NOT _509_ (
    .A(_245_),
    .Y(_246_)
  );
  NOR _510_ (
    .A(_233_),
    .B(_236_),
    .Y(_247_)
  );
  NAND _511_ (
    .A(_232_),
    .B(_237_),
    .Y(_248_)
  );
  NOR _512_ (
    .A(_234_),
    .B(_247_),
    .Y(_249_)
  );
  NAND _513_ (
    .A(_235_),
    .B(_248_),
    .Y(_250_)
  );
  NOR _514_ (
    .A(_246_),
    .B(_250_),
    .Y(_251_)
  );
  NAND _515_ (
    .A(_245_),
    .B(_249_),
    .Y(_252_)
  );
  NOR _516_ (
    .A(_245_),
    .B(_249_),
    .Y(_253_)
  );
  NOR _517_ (
    .A(_251_),
    .B(_253_),
    .Y(_117_)
  );
  NOR _518_ (
    .A(_243_),
    .B(_251_),
    .Y(_254_)
  );
  NAND _519_ (
    .A(_244_),
    .B(_252_),
    .Y(_255_)
  );
  NOR _520_ (
    .A(_102_),
    .B(_086_),
    .Y(_256_)
  );
  NAND _521_ (
    .A(_314_),
    .B(_315_),
    .Y(_257_)
  );
  NOR _522_ (
    .A(_314_),
    .B(_315_),
    .Y(_258_)
  );
  NAND _523_ (
    .A(_102_),
    .B(_086_),
    .Y(_259_)
  );
  NOR _524_ (
    .A(_256_),
    .B(_258_),
    .Y(_260_)
  );
  NAND _525_ (
    .A(_257_),
    .B(_259_),
    .Y(_261_)
  );
  NAND _526_ (
    .A(_255_),
    .B(_261_),
    .Y(_262_)
  );
  NAND _527_ (
    .A(_254_),
    .B(_260_),
    .Y(_263_)
  );
  NAND _528_ (
    .A(_262_),
    .B(_263_),
    .Y(_118_)
  );
  NOR _529_ (
    .A(_316_),
    .B(_317_),
    .Y(_264_)
  );
  NAND _530_ (
    .A(_103_),
    .B(_087_),
    .Y(_265_)
  );
  NOR _531_ (
    .A(_103_),
    .B(_087_),
    .Y(_266_)
  );
  NOR _532_ (
    .A(_264_),
    .B(_266_),
    .Y(_267_)
  );
  NOT _533_ (
    .A(_267_),
    .Y(_268_)
  );
  NOR _534_ (
    .A(_255_),
    .B(_258_),
    .Y(_269_)
  );
  NAND _535_ (
    .A(_254_),
    .B(_259_),
    .Y(_270_)
  );
  NOR _536_ (
    .A(_256_),
    .B(_269_),
    .Y(_271_)
  );
  NAND _537_ (
    .A(_257_),
    .B(_270_),
    .Y(_272_)
  );
  NOR _538_ (
    .A(_268_),
    .B(_272_),
    .Y(_273_)
  );
  NAND _539_ (
    .A(_267_),
    .B(_271_),
    .Y(_274_)
  );
  NOR _540_ (
    .A(_267_),
    .B(_271_),
    .Y(_275_)
  );
  NOR _541_ (
    .A(_273_),
    .B(_275_),
    .Y(_119_)
  );
  NOR _542_ (
    .A(_264_),
    .B(_273_),
    .Y(_276_)
  );
  NAND _543_ (
    .A(_265_),
    .B(_274_),
    .Y(_277_)
  );
  NOR _544_ (
    .A(_318_),
    .B(_319_),
    .Y(_278_)
  );
  NAND _545_ (
    .A(_104_),
    .B(_088_),
    .Y(_279_)
  );
  NOR _546_ (
    .A(_104_),
    .B(_088_),
    .Y(_280_)
  );
  NOT _547_ (
    .A(_280_),
    .Y(_281_)
  );
  NOR _548_ (
    .A(_278_),
    .B(_280_),
    .Y(_282_)
  );
  NAND _549_ (
    .A(_279_),
    .B(_281_),
    .Y(_283_)
  );
  NAND _550_ (
    .A(_277_),
    .B(_283_),
    .Y(_284_)
  );
  NAND _551_ (
    .A(_276_),
    .B(_282_),
    .Y(_285_)
  );
  NAND _552_ (
    .A(_284_),
    .B(_285_),
    .Y(_120_)
  );
  NOR _553_ (
    .A(_277_),
    .B(_278_),
    .Y(_286_)
  );
  NOR _554_ (
    .A(_280_),
    .B(_286_),
    .Y(_131_)
  );
  assign _098_ = B[0];
  assign _082_ = A[0];
  assign _130_ = ci;
  assign W[0] = _114_;
  assign _105_ = B[1];
  assign _089_ = A[1];
  assign W[1] = _121_;
  assign _106_ = B[2];
  assign _090_ = A[2];
  assign W[2] = _122_;
  assign _107_ = B[3];
  assign _091_ = A[3];
  assign W[3] = _123_;
  assign _108_ = B[4];
  assign _092_ = A[4];
  assign W[4] = _124_;
  assign _109_ = B[5];
  assign _093_ = A[5];
  assign W[5] = _125_;
  assign _110_ = B[6];
  assign _094_ = A[6];
  assign W[6] = _126_;
  assign _111_ = B[7];
  assign _095_ = A[7];
  assign W[7] = _127_;
  assign _112_ = B[8];
  assign _096_ = A[8];
  assign W[8] = _128_;
  assign _113_ = B[9];
  assign _097_ = A[9];
  assign W[9] = _129_;
  assign _099_ = B[10];
  assign _083_ = A[10];
  assign W[10] = _115_;
  assign _100_ = B[11];
  assign _084_ = A[11];
  assign W[11] = _116_;
  assign _101_ = B[12];
  assign _085_ = A[12];
  assign W[12] = _117_;
  assign _102_ = B[13];
  assign _086_ = A[13];
  assign W[13] = _118_;
  assign _103_ = B[14];
  assign _087_ = A[14];
  assign W[14] = _119_;
  assign _104_ = B[15];
  assign _088_ = A[15];
  assign W[15] = _120_;
  assign co = _131_;
endmodule

module And16bit(A, B, W);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  input [15:0] A;
  input [15:0] B;
  output [15:0] W;
  NAND _64_ (
    .A(_16_),
    .B(_00_),
    .Y(_48_)
  );
  NOT _65_ (
    .A(_48_),
    .Y(_32_)
  );
  NAND _66_ (
    .A(_23_),
    .B(_07_),
    .Y(_49_)
  );
  NOT _67_ (
    .A(_49_),
    .Y(_39_)
  );
  NAND _68_ (
    .A(_24_),
    .B(_08_),
    .Y(_50_)
  );
  NOT _69_ (
    .A(_50_),
    .Y(_40_)
  );
  NAND _70_ (
    .A(_25_),
    .B(_09_),
    .Y(_51_)
  );
  NOT _71_ (
    .A(_51_),
    .Y(_41_)
  );
  NAND _72_ (
    .A(_26_),
    .B(_10_),
    .Y(_52_)
  );
  NOT _73_ (
    .A(_52_),
    .Y(_42_)
  );
  NAND _74_ (
    .A(_27_),
    .B(_11_),
    .Y(_53_)
  );
  NOT _75_ (
    .A(_53_),
    .Y(_43_)
  );
  NAND _76_ (
    .A(_28_),
    .B(_12_),
    .Y(_54_)
  );
  NOT _77_ (
    .A(_54_),
    .Y(_44_)
  );
  NAND _78_ (
    .A(_29_),
    .B(_13_),
    .Y(_55_)
  );
  NOT _79_ (
    .A(_55_),
    .Y(_45_)
  );
  NAND _80_ (
    .A(_30_),
    .B(_14_),
    .Y(_56_)
  );
  NOT _81_ (
    .A(_56_),
    .Y(_46_)
  );
  NAND _82_ (
    .A(_31_),
    .B(_15_),
    .Y(_57_)
  );
  NOT _83_ (
    .A(_57_),
    .Y(_47_)
  );
  NAND _84_ (
    .A(_17_),
    .B(_01_),
    .Y(_58_)
  );
  NOT _85_ (
    .A(_58_),
    .Y(_33_)
  );
  NAND _86_ (
    .A(_18_),
    .B(_02_),
    .Y(_59_)
  );
  NOT _87_ (
    .A(_59_),
    .Y(_34_)
  );
  NAND _88_ (
    .A(_19_),
    .B(_03_),
    .Y(_60_)
  );
  NOT _89_ (
    .A(_60_),
    .Y(_35_)
  );
  NAND _90_ (
    .A(_20_),
    .B(_04_),
    .Y(_61_)
  );
  NOT _91_ (
    .A(_61_),
    .Y(_36_)
  );
  NAND _92_ (
    .A(_21_),
    .B(_05_),
    .Y(_62_)
  );
  NOT _93_ (
    .A(_62_),
    .Y(_37_)
  );
  NAND _94_ (
    .A(_22_),
    .B(_06_),
    .Y(_63_)
  );
  NOT _95_ (
    .A(_63_),
    .Y(_38_)
  );
  assign _16_ = B[0];
  assign _00_ = A[0];
  assign W[0] = _32_;
  assign _23_ = B[1];
  assign _07_ = A[1];
  assign W[1] = _39_;
  assign _24_ = B[2];
  assign _08_ = A[2];
  assign W[2] = _40_;
  assign _25_ = B[3];
  assign _09_ = A[3];
  assign W[3] = _41_;
  assign _26_ = B[4];
  assign _10_ = A[4];
  assign W[4] = _42_;
  assign _27_ = B[5];
  assign _11_ = A[5];
  assign W[5] = _43_;
  assign _28_ = B[6];
  assign _12_ = A[6];
  assign W[6] = _44_;
  assign _29_ = B[7];
  assign _13_ = A[7];
  assign W[7] = _45_;
  assign _30_ = B[8];
  assign _14_ = A[8];
  assign W[8] = _46_;
  assign _31_ = B[9];
  assign _15_ = A[9];
  assign W[9] = _47_;
  assign _17_ = B[10];
  assign _01_ = A[10];
  assign W[10] = _33_;
  assign _18_ = B[11];
  assign _02_ = A[11];
  assign W[11] = _34_;
  assign _19_ = B[12];
  assign _03_ = A[12];
  assign W[12] = _35_;
  assign _20_ = B[13];
  assign _04_ = A[13];
  assign W[13] = _36_;
  assign _21_ = B[14];
  assign _05_ = A[14];
  assign W[14] = _37_;
  assign _22_ = B[15];
  assign _06_ = A[15];
  assign W[15] = _38_;
endmodule

module Inventer(A, W);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  input [15:0] A;
  output [15:0] W;
  NOT _32_ (
    .A(_00_),
    .Y(_16_)
  );
  NOT _33_ (
    .A(_07_),
    .Y(_23_)
  );
  NOT _34_ (
    .A(_08_),
    .Y(_24_)
  );
  NOT _35_ (
    .A(_09_),
    .Y(_25_)
  );
  NOT _36_ (
    .A(_10_),
    .Y(_26_)
  );
  NOT _37_ (
    .A(_11_),
    .Y(_27_)
  );
  NOT _38_ (
    .A(_12_),
    .Y(_28_)
  );
  NOT _39_ (
    .A(_13_),
    .Y(_29_)
  );
  NOT _40_ (
    .A(_14_),
    .Y(_30_)
  );
  NOT _41_ (
    .A(_15_),
    .Y(_31_)
  );
  NOT _42_ (
    .A(_01_),
    .Y(_17_)
  );
  NOT _43_ (
    .A(_02_),
    .Y(_18_)
  );
  NOT _44_ (
    .A(_03_),
    .Y(_19_)
  );
  NOT _45_ (
    .A(_04_),
    .Y(_20_)
  );
  NOT _46_ (
    .A(_05_),
    .Y(_21_)
  );
  NOT _47_ (
    .A(_06_),
    .Y(_22_)
  );
  assign _00_ = A[0];
  assign W[0] = _16_;
  assign _07_ = A[1];
  assign W[1] = _23_;
  assign _08_ = A[2];
  assign W[2] = _24_;
  assign _09_ = A[3];
  assign W[3] = _25_;
  assign _10_ = A[4];
  assign W[4] = _26_;
  assign _11_ = A[5];
  assign W[5] = _27_;
  assign _12_ = A[6];
  assign W[6] = _28_;
  assign _13_ = A[7];
  assign W[7] = _29_;
  assign _14_ = A[8];
  assign W[8] = _30_;
  assign _15_ = A[9];
  assign W[9] = _31_;
  assign _01_ = A[10];
  assign W[10] = _17_;
  assign _02_ = A[11];
  assign W[11] = _18_;
  assign _03_ = A[12];
  assign W[12] = _19_;
  assign _04_ = A[13];
  assign W[13] = _20_;
  assign _05_ = A[14];
  assign W[14] = _21_;
  assign _06_ = A[15];
  assign W[15] = _22_;
endmodule

module Mux4(A1, A2, A3, A4, select, W);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  wire _257_;
  wire _258_;
  wire _259_;
  wire _260_;
  wire _261_;
  wire _262_;
  wire _263_;
  wire _264_;
  wire _265_;
  wire _266_;
  wire _267_;
  input [15:0] A1;
  input [15:0] A2;
  input [15:0] A3;
  input [15:0] A4;
  output [15:0] W;
  input [1:0] select;
  NOT _268_ (
    .A(_267_),
    .Y(_250_)
  );
  NOT _269_ (
    .A(_083_),
    .Y(_251_)
  );
  NOT _270_ (
    .A(_051_),
    .Y(_252_)
  );
  NOT _271_ (
    .A(_090_),
    .Y(_253_)
  );
  NOT _272_ (
    .A(_058_),
    .Y(_254_)
  );
  NOT _273_ (
    .A(_091_),
    .Y(_255_)
  );
  NOT _274_ (
    .A(_059_),
    .Y(_256_)
  );
  NOT _275_ (
    .A(_092_),
    .Y(_257_)
  );
  NOT _276_ (
    .A(_060_),
    .Y(_258_)
  );
  NOT _277_ (
    .A(_093_),
    .Y(_259_)
  );
  NOT _278_ (
    .A(_061_),
    .Y(_260_)
  );
  NOT _279_ (
    .A(_094_),
    .Y(_261_)
  );
  NOT _280_ (
    .A(_062_),
    .Y(_262_)
  );
  NOT _281_ (
    .A(_095_),
    .Y(_263_)
  );
  NOT _282_ (
    .A(_063_),
    .Y(_264_)
  );
  NOT _283_ (
    .A(_096_),
    .Y(_265_)
  );
  NOT _284_ (
    .A(_064_),
    .Y(_115_)
  );
  NOT _285_ (
    .A(_097_),
    .Y(_116_)
  );
  NOT _286_ (
    .A(_065_),
    .Y(_117_)
  );
  NOT _287_ (
    .A(_098_),
    .Y(_118_)
  );
  NOT _288_ (
    .A(_066_),
    .Y(_119_)
  );
  NOT _289_ (
    .A(_084_),
    .Y(_120_)
  );
  NOT _290_ (
    .A(_052_),
    .Y(_121_)
  );
  NOT _291_ (
    .A(_085_),
    .Y(_122_)
  );
  NOT _292_ (
    .A(_053_),
    .Y(_123_)
  );
  NOT _293_ (
    .A(_086_),
    .Y(_124_)
  );
  NOT _294_ (
    .A(_054_),
    .Y(_125_)
  );
  NOT _295_ (
    .A(_087_),
    .Y(_126_)
  );
  NOT _296_ (
    .A(_055_),
    .Y(_127_)
  );
  NOT _297_ (
    .A(_088_),
    .Y(_128_)
  );
  NOT _298_ (
    .A(_056_),
    .Y(_129_)
  );
  NOT _299_ (
    .A(_089_),
    .Y(_130_)
  );
  NOT _300_ (
    .A(_057_),
    .Y(_131_)
  );
  NAND _301_ (
    .A(_249_),
    .B(_250_),
    .Y(_132_)
  );
  NOR _302_ (
    .A(_035_),
    .B(_132_),
    .Y(_133_)
  );
  NAND _303_ (
    .A(_266_),
    .B(_250_),
    .Y(_134_)
  );
  NOR _304_ (
    .A(_266_),
    .B(_250_),
    .Y(_135_)
  );
  NAND _305_ (
    .A(_249_),
    .B(_267_),
    .Y(_136_)
  );
  NAND _306_ (
    .A(_134_),
    .B(_136_),
    .Y(_137_)
  );
  NOR _307_ (
    .A(_251_),
    .B(_137_),
    .Y(_138_)
  );
  NAND _308_ (
    .A(_067_),
    .B(_135_),
    .Y(_139_)
  );
  NAND _309_ (
    .A(_266_),
    .B(_252_),
    .Y(_140_)
  );
  NAND _310_ (
    .A(_250_),
    .B(_140_),
    .Y(_141_)
  );
  NAND _311_ (
    .A(_139_),
    .B(_141_),
    .Y(_142_)
  );
  NOR _312_ (
    .A(_138_),
    .B(_142_),
    .Y(_143_)
  );
  NOR _313_ (
    .A(_133_),
    .B(_143_),
    .Y(_099_)
  );
  NOR _314_ (
    .A(_042_),
    .B(_132_),
    .Y(_144_)
  );
  NOR _315_ (
    .A(_253_),
    .B(_137_),
    .Y(_145_)
  );
  NAND _316_ (
    .A(_074_),
    .B(_135_),
    .Y(_146_)
  );
  NAND _317_ (
    .A(_266_),
    .B(_254_),
    .Y(_147_)
  );
  NAND _318_ (
    .A(_250_),
    .B(_147_),
    .Y(_148_)
  );
  NAND _319_ (
    .A(_146_),
    .B(_148_),
    .Y(_149_)
  );
  NOR _320_ (
    .A(_145_),
    .B(_149_),
    .Y(_150_)
  );
  NOR _321_ (
    .A(_144_),
    .B(_150_),
    .Y(_106_)
  );
  NOR _322_ (
    .A(_043_),
    .B(_132_),
    .Y(_151_)
  );
  NOR _323_ (
    .A(_255_),
    .B(_137_),
    .Y(_152_)
  );
  NAND _324_ (
    .A(_075_),
    .B(_135_),
    .Y(_153_)
  );
  NAND _325_ (
    .A(_266_),
    .B(_256_),
    .Y(_154_)
  );
  NAND _326_ (
    .A(_250_),
    .B(_154_),
    .Y(_155_)
  );
  NAND _327_ (
    .A(_153_),
    .B(_155_),
    .Y(_156_)
  );
  NOR _328_ (
    .A(_152_),
    .B(_156_),
    .Y(_157_)
  );
  NOR _329_ (
    .A(_151_),
    .B(_157_),
    .Y(_107_)
  );
  NOR _330_ (
    .A(_044_),
    .B(_132_),
    .Y(_158_)
  );
  NOR _331_ (
    .A(_257_),
    .B(_137_),
    .Y(_159_)
  );
  NAND _332_ (
    .A(_076_),
    .B(_135_),
    .Y(_160_)
  );
  NAND _333_ (
    .A(_266_),
    .B(_258_),
    .Y(_161_)
  );
  NAND _334_ (
    .A(_250_),
    .B(_161_),
    .Y(_162_)
  );
  NAND _335_ (
    .A(_160_),
    .B(_162_),
    .Y(_163_)
  );
  NOR _336_ (
    .A(_159_),
    .B(_163_),
    .Y(_164_)
  );
  NOR _337_ (
    .A(_158_),
    .B(_164_),
    .Y(_108_)
  );
  NOR _338_ (
    .A(_045_),
    .B(_132_),
    .Y(_165_)
  );
  NOR _339_ (
    .A(_259_),
    .B(_137_),
    .Y(_166_)
  );
  NAND _340_ (
    .A(_077_),
    .B(_135_),
    .Y(_167_)
  );
  NAND _341_ (
    .A(_266_),
    .B(_260_),
    .Y(_168_)
  );
  NAND _342_ (
    .A(_250_),
    .B(_168_),
    .Y(_169_)
  );
  NAND _343_ (
    .A(_167_),
    .B(_169_),
    .Y(_170_)
  );
  NOR _344_ (
    .A(_166_),
    .B(_170_),
    .Y(_171_)
  );
  NOR _345_ (
    .A(_165_),
    .B(_171_),
    .Y(_109_)
  );
  NOR _346_ (
    .A(_046_),
    .B(_132_),
    .Y(_172_)
  );
  NOR _347_ (
    .A(_261_),
    .B(_137_),
    .Y(_173_)
  );
  NAND _348_ (
    .A(_078_),
    .B(_135_),
    .Y(_174_)
  );
  NAND _349_ (
    .A(_266_),
    .B(_262_),
    .Y(_175_)
  );
  NAND _350_ (
    .A(_250_),
    .B(_175_),
    .Y(_176_)
  );
  NAND _351_ (
    .A(_174_),
    .B(_176_),
    .Y(_177_)
  );
  NOR _352_ (
    .A(_173_),
    .B(_177_),
    .Y(_178_)
  );
  NOR _353_ (
    .A(_172_),
    .B(_178_),
    .Y(_110_)
  );
  NOR _354_ (
    .A(_047_),
    .B(_132_),
    .Y(_179_)
  );
  NOR _355_ (
    .A(_263_),
    .B(_137_),
    .Y(_180_)
  );
  NAND _356_ (
    .A(_079_),
    .B(_135_),
    .Y(_181_)
  );
  NAND _357_ (
    .A(_266_),
    .B(_264_),
    .Y(_182_)
  );
  NAND _358_ (
    .A(_250_),
    .B(_182_),
    .Y(_183_)
  );
  NAND _359_ (
    .A(_181_),
    .B(_183_),
    .Y(_184_)
  );
  NOR _360_ (
    .A(_180_),
    .B(_184_),
    .Y(_185_)
  );
  NOR _361_ (
    .A(_179_),
    .B(_185_),
    .Y(_111_)
  );
  NOR _362_ (
    .A(_048_),
    .B(_132_),
    .Y(_186_)
  );
  NOR _363_ (
    .A(_265_),
    .B(_137_),
    .Y(_187_)
  );
  NAND _364_ (
    .A(_080_),
    .B(_135_),
    .Y(_188_)
  );
  NAND _365_ (
    .A(_266_),
    .B(_115_),
    .Y(_189_)
  );
  NAND _366_ (
    .A(_250_),
    .B(_189_),
    .Y(_190_)
  );
  NAND _367_ (
    .A(_188_),
    .B(_190_),
    .Y(_191_)
  );
  NOR _368_ (
    .A(_187_),
    .B(_191_),
    .Y(_192_)
  );
  NOR _369_ (
    .A(_186_),
    .B(_192_),
    .Y(_112_)
  );
  NOR _370_ (
    .A(_049_),
    .B(_132_),
    .Y(_193_)
  );
  NOR _371_ (
    .A(_116_),
    .B(_137_),
    .Y(_194_)
  );
  NAND _372_ (
    .A(_081_),
    .B(_135_),
    .Y(_195_)
  );
  NAND _373_ (
    .A(_266_),
    .B(_117_),
    .Y(_196_)
  );
  NAND _374_ (
    .A(_250_),
    .B(_196_),
    .Y(_197_)
  );
  NAND _375_ (
    .A(_195_),
    .B(_197_),
    .Y(_198_)
  );
  NOR _376_ (
    .A(_194_),
    .B(_198_),
    .Y(_199_)
  );
  NOR _377_ (
    .A(_193_),
    .B(_199_),
    .Y(_113_)
  );
  NOR _378_ (
    .A(_050_),
    .B(_132_),
    .Y(_200_)
  );
  NOR _379_ (
    .A(_118_),
    .B(_137_),
    .Y(_201_)
  );
  NAND _380_ (
    .A(_082_),
    .B(_135_),
    .Y(_202_)
  );
  NAND _381_ (
    .A(_266_),
    .B(_119_),
    .Y(_203_)
  );
  NAND _382_ (
    .A(_250_),
    .B(_203_),
    .Y(_204_)
  );
  NAND _383_ (
    .A(_202_),
    .B(_204_),
    .Y(_205_)
  );
  NOR _384_ (
    .A(_201_),
    .B(_205_),
    .Y(_206_)
  );
  NOR _385_ (
    .A(_200_),
    .B(_206_),
    .Y(_114_)
  );
  NOR _386_ (
    .A(_036_),
    .B(_132_),
    .Y(_207_)
  );
  NOR _387_ (
    .A(_120_),
    .B(_137_),
    .Y(_208_)
  );
  NAND _388_ (
    .A(_068_),
    .B(_135_),
    .Y(_209_)
  );
  NAND _389_ (
    .A(_266_),
    .B(_121_),
    .Y(_210_)
  );
  NAND _390_ (
    .A(_250_),
    .B(_210_),
    .Y(_211_)
  );
  NAND _391_ (
    .A(_209_),
    .B(_211_),
    .Y(_212_)
  );
  NOR _392_ (
    .A(_208_),
    .B(_212_),
    .Y(_213_)
  );
  NOR _393_ (
    .A(_207_),
    .B(_213_),
    .Y(_100_)
  );
  NOR _394_ (
    .A(_037_),
    .B(_132_),
    .Y(_214_)
  );
  NOR _395_ (
    .A(_122_),
    .B(_137_),
    .Y(_215_)
  );
  NAND _396_ (
    .A(_069_),
    .B(_135_),
    .Y(_216_)
  );
  NAND _397_ (
    .A(_266_),
    .B(_123_),
    .Y(_217_)
  );
  NAND _398_ (
    .A(_250_),
    .B(_217_),
    .Y(_218_)
  );
  NAND _399_ (
    .A(_216_),
    .B(_218_),
    .Y(_219_)
  );
  NOR _400_ (
    .A(_215_),
    .B(_219_),
    .Y(_220_)
  );
  NOR _401_ (
    .A(_214_),
    .B(_220_),
    .Y(_101_)
  );
  NOR _402_ (
    .A(_038_),
    .B(_132_),
    .Y(_221_)
  );
  NOR _403_ (
    .A(_124_),
    .B(_137_),
    .Y(_222_)
  );
  NAND _404_ (
    .A(_070_),
    .B(_135_),
    .Y(_223_)
  );
  NAND _405_ (
    .A(_266_),
    .B(_125_),
    .Y(_224_)
  );
  NAND _406_ (
    .A(_250_),
    .B(_224_),
    .Y(_225_)
  );
  NAND _407_ (
    .A(_223_),
    .B(_225_),
    .Y(_226_)
  );
  NOR _408_ (
    .A(_222_),
    .B(_226_),
    .Y(_227_)
  );
  NOR _409_ (
    .A(_221_),
    .B(_227_),
    .Y(_102_)
  );
  NOR _410_ (
    .A(_039_),
    .B(_132_),
    .Y(_228_)
  );
  NOR _411_ (
    .A(_126_),
    .B(_137_),
    .Y(_229_)
  );
  NAND _412_ (
    .A(_071_),
    .B(_135_),
    .Y(_230_)
  );
  NAND _413_ (
    .A(_266_),
    .B(_127_),
    .Y(_231_)
  );
  NAND _414_ (
    .A(_250_),
    .B(_231_),
    .Y(_232_)
  );
  NAND _415_ (
    .A(_230_),
    .B(_232_),
    .Y(_233_)
  );
  NOR _416_ (
    .A(_229_),
    .B(_233_),
    .Y(_234_)
  );
  NOR _417_ (
    .A(_228_),
    .B(_234_),
    .Y(_103_)
  );
  NOR _418_ (
    .A(_040_),
    .B(_132_),
    .Y(_235_)
  );
  NOR _419_ (
    .A(_128_),
    .B(_137_),
    .Y(_236_)
  );
  NAND _420_ (
    .A(_072_),
    .B(_135_),
    .Y(_237_)
  );
  NAND _421_ (
    .A(_266_),
    .B(_129_),
    .Y(_238_)
  );
  NAND _422_ (
    .A(_250_),
    .B(_238_),
    .Y(_239_)
  );
  NAND _423_ (
    .A(_237_),
    .B(_239_),
    .Y(_240_)
  );
  NOR _424_ (
    .A(_236_),
    .B(_240_),
    .Y(_241_)
  );
  NOR _425_ (
    .A(_235_),
    .B(_241_),
    .Y(_104_)
  );
  NOR _426_ (
    .A(_041_),
    .B(_132_),
    .Y(_242_)
  );
  NOR _427_ (
    .A(_130_),
    .B(_137_),
    .Y(_243_)
  );
  NAND _428_ (
    .A(_073_),
    .B(_135_),
    .Y(_244_)
  );
  NAND _429_ (
    .A(_266_),
    .B(_131_),
    .Y(_245_)
  );
  NAND _430_ (
    .A(_250_),
    .B(_245_),
    .Y(_246_)
  );
  NAND _431_ (
    .A(_244_),
    .B(_246_),
    .Y(_247_)
  );
  NOR _432_ (
    .A(_243_),
    .B(_247_),
    .Y(_248_)
  );
  NOR _433_ (
    .A(_242_),
    .B(_248_),
    .Y(_105_)
  );
  NOT _434_ (
    .A(_266_),
    .Y(_249_)
  );
  assign _266_ = select[0];
  assign _267_ = select[1];
  assign _067_ = A3[0];
  assign _083_ = A4[0];
  assign _051_ = A2[0];
  assign _035_ = A1[0];
  assign W[0] = _099_;
  assign _074_ = A3[1];
  assign _090_ = A4[1];
  assign _058_ = A2[1];
  assign _042_ = A1[1];
  assign W[1] = _106_;
  assign _075_ = A3[2];
  assign _091_ = A4[2];
  assign _059_ = A2[2];
  assign _043_ = A1[2];
  assign W[2] = _107_;
  assign _076_ = A3[3];
  assign _092_ = A4[3];
  assign _060_ = A2[3];
  assign _044_ = A1[3];
  assign W[3] = _108_;
  assign _077_ = A3[4];
  assign _093_ = A4[4];
  assign _061_ = A2[4];
  assign _045_ = A1[4];
  assign W[4] = _109_;
  assign _078_ = A3[5];
  assign _094_ = A4[5];
  assign _062_ = A2[5];
  assign _046_ = A1[5];
  assign W[5] = _110_;
  assign _079_ = A3[6];
  assign _095_ = A4[6];
  assign _063_ = A2[6];
  assign _047_ = A1[6];
  assign W[6] = _111_;
  assign _080_ = A3[7];
  assign _096_ = A4[7];
  assign _064_ = A2[7];
  assign _048_ = A1[7];
  assign W[7] = _112_;
  assign _081_ = A3[8];
  assign _097_ = A4[8];
  assign _065_ = A2[8];
  assign _049_ = A1[8];
  assign W[8] = _113_;
  assign _082_ = A3[9];
  assign _098_ = A4[9];
  assign _066_ = A2[9];
  assign _050_ = A1[9];
  assign W[9] = _114_;
  assign _068_ = A3[10];
  assign _084_ = A4[10];
  assign _052_ = A2[10];
  assign _036_ = A1[10];
  assign W[10] = _100_;
  assign _069_ = A3[11];
  assign _085_ = A4[11];
  assign _053_ = A2[11];
  assign _037_ = A1[11];
  assign W[11] = _101_;
  assign _070_ = A3[12];
  assign _086_ = A4[12];
  assign _054_ = A2[12];
  assign _038_ = A1[12];
  assign W[12] = _102_;
  assign _071_ = A3[13];
  assign _087_ = A4[13];
  assign _055_ = A2[13];
  assign _039_ = A1[13];
  assign W[13] = _103_;
  assign _072_ = A3[14];
  assign _088_ = A4[14];
  assign _056_ = A2[14];
  assign _040_ = A1[14];
  assign W[14] = _104_;
  assign _073_ = A3[15];
  assign _089_ = A4[15];
  assign _057_ = A2[15];
  assign _041_ = A1[15];
  assign W[15] = _105_;
endmodule

module Or16bit(A, B, W);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire _53_;
  wire _54_;
  wire _55_;
  wire _56_;
  wire _57_;
  wire _58_;
  wire _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  input [15:0] A;
  input [15:0] B;
  output [15:0] W;
  NOR _64_ (
    .A(_16_),
    .B(_00_),
    .Y(_48_)
  );
  NOT _65_ (
    .A(_48_),
    .Y(_32_)
  );
  NOR _66_ (
    .A(_23_),
    .B(_07_),
    .Y(_49_)
  );
  NOT _67_ (
    .A(_49_),
    .Y(_39_)
  );
  NOR _68_ (
    .A(_24_),
    .B(_08_),
    .Y(_50_)
  );
  NOT _69_ (
    .A(_50_),
    .Y(_40_)
  );
  NOR _70_ (
    .A(_25_),
    .B(_09_),
    .Y(_51_)
  );
  NOT _71_ (
    .A(_51_),
    .Y(_41_)
  );
  NOR _72_ (
    .A(_26_),
    .B(_10_),
    .Y(_52_)
  );
  NOT _73_ (
    .A(_52_),
    .Y(_42_)
  );
  NOR _74_ (
    .A(_27_),
    .B(_11_),
    .Y(_53_)
  );
  NOT _75_ (
    .A(_53_),
    .Y(_43_)
  );
  NOR _76_ (
    .A(_28_),
    .B(_12_),
    .Y(_54_)
  );
  NOT _77_ (
    .A(_54_),
    .Y(_44_)
  );
  NOR _78_ (
    .A(_29_),
    .B(_13_),
    .Y(_55_)
  );
  NOT _79_ (
    .A(_55_),
    .Y(_45_)
  );
  NOR _80_ (
    .A(_30_),
    .B(_14_),
    .Y(_56_)
  );
  NOT _81_ (
    .A(_56_),
    .Y(_46_)
  );
  NOR _82_ (
    .A(_31_),
    .B(_15_),
    .Y(_57_)
  );
  NOT _83_ (
    .A(_57_),
    .Y(_47_)
  );
  NOR _84_ (
    .A(_17_),
    .B(_01_),
    .Y(_58_)
  );
  NOT _85_ (
    .A(_58_),
    .Y(_33_)
  );
  NOR _86_ (
    .A(_18_),
    .B(_02_),
    .Y(_59_)
  );
  NOT _87_ (
    .A(_59_),
    .Y(_34_)
  );
  NOR _88_ (
    .A(_19_),
    .B(_03_),
    .Y(_60_)
  );
  NOT _89_ (
    .A(_60_),
    .Y(_35_)
  );
  NOR _90_ (
    .A(_20_),
    .B(_04_),
    .Y(_61_)
  );
  NOT _91_ (
    .A(_61_),
    .Y(_36_)
  );
  NOR _92_ (
    .A(_21_),
    .B(_05_),
    .Y(_62_)
  );
  NOT _93_ (
    .A(_62_),
    .Y(_37_)
  );
  NOR _94_ (
    .A(_22_),
    .B(_06_),
    .Y(_63_)
  );
  NOT _95_ (
    .A(_63_),
    .Y(_38_)
  );
  assign _16_ = B[0];
  assign _00_ = A[0];
  assign W[0] = _32_;
  assign _23_ = B[1];
  assign _07_ = A[1];
  assign W[1] = _39_;
  assign _24_ = B[2];
  assign _08_ = A[2];
  assign W[2] = _40_;
  assign _25_ = B[3];
  assign _09_ = A[3];
  assign W[3] = _41_;
  assign _26_ = B[4];
  assign _10_ = A[4];
  assign W[4] = _42_;
  assign _27_ = B[5];
  assign _11_ = A[5];
  assign W[5] = _43_;
  assign _28_ = B[6];
  assign _12_ = A[6];
  assign W[6] = _44_;
  assign _29_ = B[7];
  assign _13_ = A[7];
  assign W[7] = _45_;
  assign _30_ = B[8];
  assign _14_ = A[8];
  assign W[8] = _46_;
  assign _31_ = B[9];
  assign _15_ = A[9];
  assign W[9] = _47_;
  assign _17_ = B[10];
  assign _01_ = A[10];
  assign W[10] = _33_;
  assign _18_ = B[11];
  assign _02_ = A[11];
  assign W[11] = _34_;
  assign _19_ = B[12];
  assign _03_ = A[12];
  assign W[12] = _35_;
  assign _20_ = B[13];
  assign _04_ = A[13];
  assign W[13] = _36_;
  assign _21_ = B[14];
  assign _05_ = A[14];
  assign W[14] = _37_;
  assign _22_ = B[15];
  assign _06_ = A[15];
  assign W[15] = _38_;
endmodule

module Orbits(A, W);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire _15_;
  wire _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  input [15:0] A;
  output W;
  NOR _45_ (
    .A(_02_),
    .B(_14_),
    .Y(_17_)
  );
  NOR _46_ (
    .A(_05_),
    .B(_04_),
    .Y(_18_)
  );
  NAND _47_ (
    .A(_17_),
    .B(_18_),
    .Y(_19_)
  );
  NOR _48_ (
    .A(_08_),
    .B(_07_),
    .Y(_20_)
  );
  NOR _49_ (
    .A(_13_),
    .B(_10_),
    .Y(_21_)
  );
  NAND _50_ (
    .A(_20_),
    .B(_21_),
    .Y(_22_)
  );
  NOR _51_ (
    .A(_19_),
    .B(_22_),
    .Y(_23_)
  );
  NOR _52_ (
    .A(_01_),
    .B(_15_),
    .Y(_24_)
  );
  NOR _53_ (
    .A(_06_),
    .B(_03_),
    .Y(_25_)
  );
  NAND _54_ (
    .A(_24_),
    .B(_25_),
    .Y(_26_)
  );
  NOR _55_ (
    .A(_09_),
    .B(_00_),
    .Y(_27_)
  );
  NOR _56_ (
    .A(_12_),
    .B(_11_),
    .Y(_28_)
  );
  NAND _57_ (
    .A(_27_),
    .B(_28_),
    .Y(_29_)
  );
  NOR _58_ (
    .A(_26_),
    .B(_29_),
    .Y(_30_)
  );
  NAND _59_ (
    .A(_23_),
    .B(_30_),
    .Y(_16_)
  );
  assign _05_ = A[14];
  assign _06_ = A[15];
  assign _03_ = A[12];
  assign _04_ = A[13];
  assign _01_ = A[10];
  assign _02_ = A[11];
  assign _14_ = A[8];
  assign _15_ = A[9];
  assign _12_ = A[6];
  assign _13_ = A[7];
  assign _10_ = A[4];
  assign _11_ = A[5];
  assign _08_ = A[2];
  assign _09_ = A[3];
  assign _00_ = A[0];
  assign _07_ = A[1];
  assign W = _16_;
endmodule

module Q2_yosys(inM, inN, inC, opc, outF, zer, neg);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire _12_;
  wire [14:0] _13_;
  wire co;
  input inC;
  input [15:0] inM;
  input [15:0] inN;
  output neg;
  input [2:0] opc;
  output [15:0] outF;
  wire w3;
  wire w4;
  wire w5;
  wire w6;
  wire wAdd;
  wire [15:0] wAnd;
  wire [15:0] wInv;
  wire [15:0] wMux;
  wire [15:0] wOr;
  wire [15:0] wShif1;
  wire [15:0] wShif2;
  output zer;
  NOT _14_ (
    .A(_09_),
    .Y(_11_)
  );
  NOT _15_ (
    .A(_04_),
    .Y(_00_)
  );
  NOT _16_ (
    .A(_06_),
    .Y(_01_)
  );
  NOR _17_ (
    .A(_05_),
    .B(_04_),
    .Y(_02_)
  );
  NOT _18_ (
    .A(_02_),
    .Y(_03_)
  );
  NOR _19_ (
    .A(_06_),
    .B(_03_),
    .Y(_10_)
  );
  NOR _20_ (
    .A(_01_),
    .B(_02_),
    .Y(_07_)
  );
  NOR _21_ (
    .A(_00_),
    .B(_06_),
    .Y(_08_)
  );
  Adder A1 (
    .A(inM),
    .B(wMux),
    .W({ _13_, co }),
    .ci(w6),
    .co(wAdd)
  );
  Inventer G1 (
    .A(inM),
    .W(wInv)
  );
  Or16bit G2 (
    .A(inM),
    .B(inN),
    .W(wOr)
  );
  And16bit G3 (
    .A(inM),
    .B(inN),
    .W(wAnd)
  );
  Orbits G4 (
    .A(outF),
    .W(w5)
  );
  Mux4 M1 (
    .A1({ 15'h0000, wAdd }),
    .A2(wAnd),
    .A3(wOr),
    .A4(wInv),
    .W(outF),
    .select({ w3, w4 })
  );
  Mux4 M2 (
    .A1(inN),
    .A2(wShif1),
    .A3(16'h0001),
    .A4(wShif2),
    .W(wMux),
    .select(opc[1:0])
  );
  Shifter2bit1 S1 (
    .A(inN),
    .W(wShif1)
  );
  Shifter2bit1 S2 (
    .A(inM),
    .W(wShif2)
  );
  assign neg = outF[15];
  assign _09_ = w5;
  assign zer = _11_;
  assign _05_ = opc[1];
  assign _04_ = opc[0];
  assign _06_ = opc[2];
  assign w6 = _10_;
  assign w3 = _07_;
  assign w4 = _08_;
endmodule

module Shifter2bit1(A, W);
  input [15:0] A;
  output [15:0] W;
  assign W = { A[15], A[15:1] };
endmodule
